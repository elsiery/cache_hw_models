/*
MIT License

Copyright (c) 2024 Elsie Rezinold Y

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.
*/
module fw_associative #(
    parameter ADDRESS_WIDTH =64,
    parameter WRITE_DATA=64,
    parameter BLOCK_SIZE_BYTE=64,
    parameter BLOCK_SIZE_BITS=6,
    parameter BLOCK_NUMBER_BITS=10,
    parameter SET_BITS = 2,
    parameter BLOCK_NUMBER = 256,
    parameter CACHE_SIZE=64*1024
)(
clk,
rst_n,
i_cpu_valid,
i_cpu_rd_wr,
i_cpu_address,
i_cpu_wr_data,
o_cpu_rd_data,
o_cpu_busy,

o_mem_rd_en,
o_mem_rd_address,
o_mem_wr_en,
o_mem_wr_address,
o_mem_wr_data,
i_mem_rd_data,
i_mem_rd_valid
);

input clk;
input rst_n;
localparam TAG_WIDTH = ADDRESS_WIDTH-(BLOCK_NUMBER_BITS - SET_BITS)-BLOCK_SIZE_BITS;
localparam BLOCK_ADDRESS_HIGH = ADDRESS_WIDTH-TAG_WIDTH-1;
localparam BLOCK_ADDRESS_LOW = BLOCK_SIZE_BITS; 
localparam TAG_HIGH = ADDRESS_WIDTH-1;
localparam TAG_LOW = BLOCK_ADDRESS_HIGH +1; 
input i_cpu_valid;
input i_cpu_rd_wr;
input [ADDRESS_WIDTH-1:0] i_cpu_address;

input [WRITE_DATA*8-1:0] i_cpu_wr_data;
output reg [WRITE_DATA*8-1:0] o_cpu_rd_data;
output reg o_cpu_busy;
output o_mem_rd_en;
output [ADDRESS_WIDTH-1:0] o_mem_rd_address;
output reg o_mem_wr_en;
output reg [ADDRESS_WIDTH-1:0] o_mem_wr_address;
output reg [WRITE_DATA*8-1:0] o_mem_wr_data;
input [WRITE_DATA*8-1:0] i_mem_rd_data;
input i_mem_rd_valid;
localparam CACHE_ACCESS=0,MISS=1;

reg [BLOCK_SIZE_BYTE*8-1:0] cache_block_1 [0:BLOCK_NUMBER-1];
reg valid_bit_1 [0:BLOCK_NUMBER-1];
reg dirty_bit_1 [0:BLOCK_NUMBER-1];
reg [TAG_WIDTH-1:0] tag_address_1[0:BLOCK_NUMBER-1];
reg [1:0] lru_counter_1 [0:BLOCK_NUMBER-1];

reg [BLOCK_SIZE_BYTE*8-1:0] cache_block_2 [0:BLOCK_NUMBER-1];
reg valid_bit_2 [0:BLOCK_NUMBER-1];
reg dirty_bit_2 [0:BLOCK_NUMBER-1];
reg [TAG_WIDTH-1:0] tag_address_2[0:BLOCK_NUMBER-1];
reg [1:0] lru_counter_2 [0:BLOCK_NUMBER-1];

reg [BLOCK_SIZE_BYTE*8-1:0] cache_block_3 [0:BLOCK_NUMBER-1];
reg valid_bit_3 [0:BLOCK_NUMBER-1];
reg dirty_bit_3 [0:BLOCK_NUMBER-1];
reg [TAG_WIDTH-1:0] tag_address_3[0:BLOCK_NUMBER-1];
reg [1:0] lru_counter_3 [0:BLOCK_NUMBER-1];

reg [BLOCK_SIZE_BYTE*8-1:0] cache_block_4 [0:BLOCK_NUMBER-1];
reg valid_bit_4 [0:BLOCK_NUMBER-1];
reg dirty_bit_4 [0:BLOCK_NUMBER-1];
reg [TAG_WIDTH-1:0] tag_address_4[0:BLOCK_NUMBER-1];
reg [1:0] lru_counter_4 [0:BLOCK_NUMBER-1];







reg cs,ns;
wire miss;
reg handled; 

assign miss = i_cpu_valid && ((i_cpu_address[TAG_HIGH:TAG_LOW]!=tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) || !valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])
                                          && ((i_cpu_address[TAG_HIGH:TAG_LOW]!=tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) || !valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])
                                          && ((i_cpu_address[TAG_HIGH:TAG_LOW]!=tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) || !valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])
                                          && ((i_cpu_address[TAG_HIGH:TAG_LOW]!=tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) || !valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]);


//assign hit  = i_cpu_valid&((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])&valid_bit[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]); 

always@(posedge clk or negedge rst_n) begin
    if(!rst_n)
        cs <= 0;
    else    
        cs <= ns;
end



always @(*) begin
    ns = 0;
    case(cs)
    CACHE_ACCESS: begin 
        if(miss) begin
            ns = MISS;
        end
    end
    MISS: begin
        if(handled) begin
            ns = CACHE_ACCESS;
        end 
        else begin
            ns = MISS;
        end
    end
    endcase
end
assign o_mem_rd_en = miss;
assign o_mem_rd_address = i_cpu_address;
always@(posedge clk or negedge rst_n) begin
    if(rst_n) begin
        case(cs)
        CACHE_ACCESS: begin
            handled <=0;
            o_mem_wr_en <=0;
            if(i_cpu_valid & !i_cpu_rd_wr) begin
                if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //rd hit 
                    //BLOCK 1
                    o_cpu_rd_data                                                       <= cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    o_cpu_busy                                                          <= 0;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //rd hit 
                    //BLOCK 2
                    o_cpu_rd_data                                                       <= cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    o_cpu_busy                                                          <= 0;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //rd hit 
                    //BLOCK 3
                    o_cpu_rd_data                                                       <= cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    o_cpu_busy                                                          <= 0;
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //rd hit 
                    //BLOCK 4
                    o_cpu_rd_data                                                       <= cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    o_cpu_busy                                                          <= 0;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else begin
                    o_cpu_busy       <= 1;
                end
            end
            else if(i_cpu_valid & i_cpu_rd_wr) begin
                if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //wr hit
                    //block 1
                    cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= i_cpu_wr_data;
                    dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]    <= 1;
                    o_cpu_busy                                                          <= 0;
                    o_mem_wr_en                                                         <= 0;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //wr hit
                    //block 2
                    cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= i_cpu_wr_data;
                    dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]    <= 1;
                    o_cpu_busy                                                          <= 0;
                    o_mem_wr_en                                                         <= 0;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //wr hit
                    //block 3
                    cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= i_cpu_wr_data;
                    dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]    <= 1;
                    o_cpu_busy                                                          <= 0;
                    o_mem_wr_en                                                         <= 0;
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else if((i_cpu_address[TAG_HIGH:TAG_LOW]==tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) && valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                    //wr hit
                    //block 4
                    cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= i_cpu_wr_data;
                    dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]    <= 1;
                    o_cpu_busy                                                          <= 0;
                    o_mem_wr_en                                                         <= 0;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
                else begin
                    o_cpu_busy<=1;
                end
            end
        end
        MISS: begin
            if(!valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                if(i_mem_rd_valid) begin                
                    cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
                    handled                                                                  <=   1;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2; 
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0; 
                end
            end
            else if(!valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                if(i_mem_rd_valid) begin                
                    cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
                    handled                                                                  <=   1;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3; 
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0; 
                end
            end
            else if(!valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                if(i_mem_rd_valid) begin                
                    cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
                    handled                                                                  <=   1;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2; 
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0; 
                end
            end
            else if(!valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                if(i_mem_rd_valid) begin                
                    cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
                    handled                                                                  <=   1;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1; 
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3; 
                end
            end
            else if(lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
                if(i_mem_rd_valid) begin                
                    if(dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                        o_mem_wr_data <= cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                        o_mem_wr_address <= {tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};;
                        o_mem_wr_en <= 1;
                    end
                    cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    handled                                                                  <=   1;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                
                end
            end
            else if(lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
                if(i_mem_rd_valid) begin                
                    if(dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                        o_mem_wr_data <= cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                        o_mem_wr_address <= {tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
                        o_mem_wr_en <= 1;
                    end
                    cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    handled                                                                  <=   1;
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                
                end
            end
            else if(lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
                if(i_mem_rd_valid) begin                
                    if(dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                        o_mem_wr_data <= cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                        o_mem_wr_address <= {tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
                        o_mem_wr_en <= 1;
                    end
                    cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    handled                                                                  <=   1;
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
            end
            else if(lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
                if(i_mem_rd_valid) begin                
                    if(dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
                        o_mem_wr_data <= cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                        o_mem_wr_address <= {tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
                        o_mem_wr_en <= 1;
                    end
                    cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_mem_rd_data;
                    tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
                    dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   0;
                    handled                                                                  <=   1;
                    lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
                    lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                    lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
                end
            end
        end
        endcase
    end
    else if(!rst_n) begin
        o_cpu_rd_data<=0;
        o_cpu_busy<=0;
        o_mem_wr_address<=0;
        o_mem_wr_en<=0;
        o_mem_wr_data<=0;
        valid_bit_1[0]  <=   0;dirty_bit_1[0] <= 0;tag_address_1[0] <= 0;cache_block_1[0] <= 0;lru_counter_1[0] <= 0;valid_bit_2[0]  <=   0;dirty_bit_2[0] <= 0;tag_address_2[0] <= 0;cache_block_2[0] <= 0;lru_counter_2[0] <= 0;valid_bit_3[0]  <=   0;dirty_bit_3[0] <= 0;tag_address_3[0] <= 0;cache_block_3[0] <= 0;lru_counter_3[0] <= 0;valid_bit_4[0]  <=   0;dirty_bit_4[0] <= 0;tag_address_4[0] <= 0;cache_block_4[0] <= 0;lru_counter_4[0] <= 0;
        valid_bit_1[1]  <=   0;dirty_bit_1[1] <= 0;tag_address_1[1] <= 0;cache_block_1[1] <= 0;lru_counter_1[1] <= 0;valid_bit_2[1]  <=   0;dirty_bit_2[1] <= 0;tag_address_2[1] <= 0;cache_block_2[1] <= 0;lru_counter_2[1] <= 0;valid_bit_3[1]  <=   0;dirty_bit_3[1] <= 0;tag_address_3[1] <= 0;cache_block_3[1] <= 0;lru_counter_3[1] <= 0;valid_bit_4[1]  <=   0;dirty_bit_4[1] <= 0;tag_address_4[1] <= 0;cache_block_4[1] <= 0;lru_counter_4[1] <= 0;
        valid_bit_1[2]  <=   0;dirty_bit_1[2] <= 0;tag_address_1[2] <= 0;cache_block_1[2] <= 0;lru_counter_1[2] <= 0;valid_bit_2[2]  <=   0;dirty_bit_2[2] <= 0;tag_address_2[2] <= 0;cache_block_2[2] <= 0;lru_counter_2[2] <= 0;valid_bit_3[2]  <=   0;dirty_bit_3[2] <= 0;tag_address_3[2] <= 0;cache_block_3[2] <= 0;lru_counter_3[2] <= 0;valid_bit_4[2]  <=   0;dirty_bit_4[2] <= 0;tag_address_4[2] <= 0;cache_block_4[2] <= 0;lru_counter_4[2] <= 0;
        valid_bit_1[3]  <=   0;dirty_bit_1[3] <= 0;tag_address_1[3] <= 0;cache_block_1[3] <= 0;lru_counter_1[3] <= 0;valid_bit_2[3]  <=   0;dirty_bit_2[3] <= 0;tag_address_2[3] <= 0;cache_block_2[3] <= 0;lru_counter_2[3] <= 0;valid_bit_3[3]  <=   0;dirty_bit_3[3] <= 0;tag_address_3[3] <= 0;cache_block_3[3] <= 0;lru_counter_3[3] <= 0;valid_bit_4[3]  <=   0;dirty_bit_4[3] <= 0;tag_address_4[3] <= 0;cache_block_4[3] <= 0;lru_counter_4[3] <= 0;
        valid_bit_1[4]  <=   0;dirty_bit_1[4] <= 0;tag_address_1[4] <= 0;cache_block_1[4] <= 0;lru_counter_1[4] <= 0;valid_bit_2[4]  <=   0;dirty_bit_2[4] <= 0;tag_address_2[4] <= 0;cache_block_2[4] <= 0;lru_counter_2[4] <= 0;valid_bit_3[4]  <=   0;dirty_bit_3[4] <= 0;tag_address_3[4] <= 0;cache_block_3[4] <= 0;lru_counter_3[4] <= 0;valid_bit_4[4]  <=   0;dirty_bit_4[4] <= 0;tag_address_4[4] <= 0;cache_block_4[4] <= 0;lru_counter_4[4] <= 0;
        valid_bit_1[5]  <=   0;dirty_bit_1[5] <= 0;tag_address_1[5] <= 0;cache_block_1[5] <= 0;lru_counter_1[5] <= 0;valid_bit_2[5]  <=   0;dirty_bit_2[5] <= 0;tag_address_2[5] <= 0;cache_block_2[5] <= 0;lru_counter_2[5] <= 0;valid_bit_3[5]  <=   0;dirty_bit_3[5] <= 0;tag_address_3[5] <= 0;cache_block_3[5] <= 0;lru_counter_3[5] <= 0;valid_bit_4[5]  <=   0;dirty_bit_4[5] <= 0;tag_address_4[5] <= 0;cache_block_4[5] <= 0;lru_counter_4[5] <= 0;
        valid_bit_1[6]  <=   0;dirty_bit_1[6] <= 0;tag_address_1[6] <= 0;cache_block_1[6] <= 0;lru_counter_1[6] <= 0;valid_bit_2[6]  <=   0;dirty_bit_2[6] <= 0;tag_address_2[6] <= 0;cache_block_2[6] <= 0;lru_counter_2[6] <= 0;valid_bit_3[6]  <=   0;dirty_bit_3[6] <= 0;tag_address_3[6] <= 0;cache_block_3[6] <= 0;lru_counter_3[6] <= 0;valid_bit_4[6]  <=   0;dirty_bit_4[6] <= 0;tag_address_4[6] <= 0;cache_block_4[6] <= 0;lru_counter_4[6] <= 0;
        valid_bit_1[7]  <=   0;dirty_bit_1[7] <= 0;tag_address_1[7] <= 0;cache_block_1[7] <= 0;lru_counter_1[7] <= 0;valid_bit_2[7]  <=   0;dirty_bit_2[7] <= 0;tag_address_2[7] <= 0;cache_block_2[7] <= 0;lru_counter_2[7] <= 0;valid_bit_3[7]  <=   0;dirty_bit_3[7] <= 0;tag_address_3[7] <= 0;cache_block_3[7] <= 0;lru_counter_3[7] <= 0;valid_bit_4[7]  <=   0;dirty_bit_4[7] <= 0;tag_address_4[7] <= 0;cache_block_4[7] <= 0;lru_counter_4[7] <= 0;
        valid_bit_1[8]  <=   0;dirty_bit_1[8] <= 0;tag_address_1[8] <= 0;cache_block_1[8] <= 0;lru_counter_1[8] <= 0;valid_bit_2[8]  <=   0;dirty_bit_2[8] <= 0;tag_address_2[8] <= 0;cache_block_2[8] <= 0;lru_counter_2[8] <= 0;valid_bit_3[8]  <=   0;dirty_bit_3[8] <= 0;tag_address_3[8] <= 0;cache_block_3[8] <= 0;lru_counter_3[8] <= 0;valid_bit_4[8]  <=   0;dirty_bit_4[8] <= 0;tag_address_4[8] <= 0;cache_block_4[8] <= 0;lru_counter_4[8] <= 0;
        valid_bit_1[9]  <=   0;dirty_bit_1[9] <= 0;tag_address_1[9] <= 0;cache_block_1[9] <= 0;lru_counter_1[9] <= 0;valid_bit_2[9]  <=   0;dirty_bit_2[9] <= 0;tag_address_2[9] <= 0;cache_block_2[9] <= 0;lru_counter_2[9] <= 0;valid_bit_3[9]  <=   0;dirty_bit_3[9] <= 0;tag_address_3[9] <= 0;cache_block_3[9] <= 0;lru_counter_3[9] <= 0;valid_bit_4[9]  <=   0;dirty_bit_4[9] <= 0;tag_address_4[9] <= 0;cache_block_4[9] <= 0;lru_counter_4[9] <= 0;
        valid_bit_1[10]  <=   0;dirty_bit_1[10] <= 0;tag_address_1[10] <= 0;cache_block_1[10] <= 0;lru_counter_1[10] <= 0;valid_bit_2[10]  <=   0;dirty_bit_2[10] <= 0;tag_address_2[10] <= 0;cache_block_2[10] <= 0;lru_counter_2[10] <= 0;valid_bit_3[10]  <=   0;dirty_bit_3[10] <= 0;tag_address_3[10] <= 0;cache_block_3[10] <= 0;lru_counter_3[10] <= 0;valid_bit_4[10]  <=   0;dirty_bit_4[10] <= 0;tag_address_4[10] <= 0;cache_block_4[10] <= 0;lru_counter_4[10] <= 0;
        valid_bit_1[11]  <=   0;dirty_bit_1[11] <= 0;tag_address_1[11] <= 0;cache_block_1[11] <= 0;lru_counter_1[11] <= 0;valid_bit_2[11]  <=   0;dirty_bit_2[11] <= 0;tag_address_2[11] <= 0;cache_block_2[11] <= 0;lru_counter_2[11] <= 0;valid_bit_3[11]  <=   0;dirty_bit_3[11] <= 0;tag_address_3[11] <= 0;cache_block_3[11] <= 0;lru_counter_3[11] <= 0;valid_bit_4[11]  <=   0;dirty_bit_4[11] <= 0;tag_address_4[11] <= 0;cache_block_4[11] <= 0;lru_counter_4[11] <= 0;
        valid_bit_1[12]  <=   0;dirty_bit_1[12] <= 0;tag_address_1[12] <= 0;cache_block_1[12] <= 0;lru_counter_1[12] <= 0;valid_bit_2[12]  <=   0;dirty_bit_2[12] <= 0;tag_address_2[12] <= 0;cache_block_2[12] <= 0;lru_counter_2[12] <= 0;valid_bit_3[12]  <=   0;dirty_bit_3[12] <= 0;tag_address_3[12] <= 0;cache_block_3[12] <= 0;lru_counter_3[12] <= 0;valid_bit_4[12]  <=   0;dirty_bit_4[12] <= 0;tag_address_4[12] <= 0;cache_block_4[12] <= 0;lru_counter_4[12] <= 0;
        valid_bit_1[13]  <=   0;dirty_bit_1[13] <= 0;tag_address_1[13] <= 0;cache_block_1[13] <= 0;lru_counter_1[13] <= 0;valid_bit_2[13]  <=   0;dirty_bit_2[13] <= 0;tag_address_2[13] <= 0;cache_block_2[13] <= 0;lru_counter_2[13] <= 0;valid_bit_3[13]  <=   0;dirty_bit_3[13] <= 0;tag_address_3[13] <= 0;cache_block_3[13] <= 0;lru_counter_3[13] <= 0;valid_bit_4[13]  <=   0;dirty_bit_4[13] <= 0;tag_address_4[13] <= 0;cache_block_4[13] <= 0;lru_counter_4[13] <= 0;
        valid_bit_1[14]  <=   0;dirty_bit_1[14] <= 0;tag_address_1[14] <= 0;cache_block_1[14] <= 0;lru_counter_1[14] <= 0;valid_bit_2[14]  <=   0;dirty_bit_2[14] <= 0;tag_address_2[14] <= 0;cache_block_2[14] <= 0;lru_counter_2[14] <= 0;valid_bit_3[14]  <=   0;dirty_bit_3[14] <= 0;tag_address_3[14] <= 0;cache_block_3[14] <= 0;lru_counter_3[14] <= 0;valid_bit_4[14]  <=   0;dirty_bit_4[14] <= 0;tag_address_4[14] <= 0;cache_block_4[14] <= 0;lru_counter_4[14] <= 0;
        valid_bit_1[15]  <=   0;dirty_bit_1[15] <= 0;tag_address_1[15] <= 0;cache_block_1[15] <= 0;lru_counter_1[15] <= 0;valid_bit_2[15]  <=   0;dirty_bit_2[15] <= 0;tag_address_2[15] <= 0;cache_block_2[15] <= 0;lru_counter_2[15] <= 0;valid_bit_3[15]  <=   0;dirty_bit_3[15] <= 0;tag_address_3[15] <= 0;cache_block_3[15] <= 0;lru_counter_3[15] <= 0;valid_bit_4[15]  <=   0;dirty_bit_4[15] <= 0;tag_address_4[15] <= 0;cache_block_4[15] <= 0;lru_counter_4[15] <= 0;
        valid_bit_1[16]  <=   0;dirty_bit_1[16] <= 0;tag_address_1[16] <= 0;cache_block_1[16] <= 0;lru_counter_1[16] <= 0;valid_bit_2[16]  <=   0;dirty_bit_2[16] <= 0;tag_address_2[16] <= 0;cache_block_2[16] <= 0;lru_counter_2[16] <= 0;valid_bit_3[16]  <=   0;dirty_bit_3[16] <= 0;tag_address_3[16] <= 0;cache_block_3[16] <= 0;lru_counter_3[16] <= 0;valid_bit_4[16]  <=   0;dirty_bit_4[16] <= 0;tag_address_4[16] <= 0;cache_block_4[16] <= 0;lru_counter_4[16] <= 0;
        valid_bit_1[17]  <=   0;dirty_bit_1[17] <= 0;tag_address_1[17] <= 0;cache_block_1[17] <= 0;lru_counter_1[17] <= 0;valid_bit_2[17]  <=   0;dirty_bit_2[17] <= 0;tag_address_2[17] <= 0;cache_block_2[17] <= 0;lru_counter_2[17] <= 0;valid_bit_3[17]  <=   0;dirty_bit_3[17] <= 0;tag_address_3[17] <= 0;cache_block_3[17] <= 0;lru_counter_3[17] <= 0;valid_bit_4[17]  <=   0;dirty_bit_4[17] <= 0;tag_address_4[17] <= 0;cache_block_4[17] <= 0;lru_counter_4[17] <= 0;
        valid_bit_1[18]  <=   0;dirty_bit_1[18] <= 0;tag_address_1[18] <= 0;cache_block_1[18] <= 0;lru_counter_1[18] <= 0;valid_bit_2[18]  <=   0;dirty_bit_2[18] <= 0;tag_address_2[18] <= 0;cache_block_2[18] <= 0;lru_counter_2[18] <= 0;valid_bit_3[18]  <=   0;dirty_bit_3[18] <= 0;tag_address_3[18] <= 0;cache_block_3[18] <= 0;lru_counter_3[18] <= 0;valid_bit_4[18]  <=   0;dirty_bit_4[18] <= 0;tag_address_4[18] <= 0;cache_block_4[18] <= 0;lru_counter_4[18] <= 0;
        valid_bit_1[19]  <=   0;dirty_bit_1[19] <= 0;tag_address_1[19] <= 0;cache_block_1[19] <= 0;lru_counter_1[19] <= 0;valid_bit_2[19]  <=   0;dirty_bit_2[19] <= 0;tag_address_2[19] <= 0;cache_block_2[19] <= 0;lru_counter_2[19] <= 0;valid_bit_3[19]  <=   0;dirty_bit_3[19] <= 0;tag_address_3[19] <= 0;cache_block_3[19] <= 0;lru_counter_3[19] <= 0;valid_bit_4[19]  <=   0;dirty_bit_4[19] <= 0;tag_address_4[19] <= 0;cache_block_4[19] <= 0;lru_counter_4[19] <= 0;
        valid_bit_1[20]  <=   0;dirty_bit_1[20] <= 0;tag_address_1[20] <= 0;cache_block_1[20] <= 0;lru_counter_1[20] <= 0;valid_bit_2[20]  <=   0;dirty_bit_2[20] <= 0;tag_address_2[20] <= 0;cache_block_2[20] <= 0;lru_counter_2[20] <= 0;valid_bit_3[20]  <=   0;dirty_bit_3[20] <= 0;tag_address_3[20] <= 0;cache_block_3[20] <= 0;lru_counter_3[20] <= 0;valid_bit_4[20]  <=   0;dirty_bit_4[20] <= 0;tag_address_4[20] <= 0;cache_block_4[20] <= 0;lru_counter_4[20] <= 0;
        valid_bit_1[21]  <=   0;dirty_bit_1[21] <= 0;tag_address_1[21] <= 0;cache_block_1[21] <= 0;lru_counter_1[21] <= 0;valid_bit_2[21]  <=   0;dirty_bit_2[21] <= 0;tag_address_2[21] <= 0;cache_block_2[21] <= 0;lru_counter_2[21] <= 0;valid_bit_3[21]  <=   0;dirty_bit_3[21] <= 0;tag_address_3[21] <= 0;cache_block_3[21] <= 0;lru_counter_3[21] <= 0;valid_bit_4[21]  <=   0;dirty_bit_4[21] <= 0;tag_address_4[21] <= 0;cache_block_4[21] <= 0;lru_counter_4[21] <= 0;
        valid_bit_1[22]  <=   0;dirty_bit_1[22] <= 0;tag_address_1[22] <= 0;cache_block_1[22] <= 0;lru_counter_1[22] <= 0;valid_bit_2[22]  <=   0;dirty_bit_2[22] <= 0;tag_address_2[22] <= 0;cache_block_2[22] <= 0;lru_counter_2[22] <= 0;valid_bit_3[22]  <=   0;dirty_bit_3[22] <= 0;tag_address_3[22] <= 0;cache_block_3[22] <= 0;lru_counter_3[22] <= 0;valid_bit_4[22]  <=   0;dirty_bit_4[22] <= 0;tag_address_4[22] <= 0;cache_block_4[22] <= 0;lru_counter_4[22] <= 0;
        valid_bit_1[23]  <=   0;dirty_bit_1[23] <= 0;tag_address_1[23] <= 0;cache_block_1[23] <= 0;lru_counter_1[23] <= 0;valid_bit_2[23]  <=   0;dirty_bit_2[23] <= 0;tag_address_2[23] <= 0;cache_block_2[23] <= 0;lru_counter_2[23] <= 0;valid_bit_3[23]  <=   0;dirty_bit_3[23] <= 0;tag_address_3[23] <= 0;cache_block_3[23] <= 0;lru_counter_3[23] <= 0;valid_bit_4[23]  <=   0;dirty_bit_4[23] <= 0;tag_address_4[23] <= 0;cache_block_4[23] <= 0;lru_counter_4[23] <= 0;
        valid_bit_1[24]  <=   0;dirty_bit_1[24] <= 0;tag_address_1[24] <= 0;cache_block_1[24] <= 0;lru_counter_1[24] <= 0;valid_bit_2[24]  <=   0;dirty_bit_2[24] <= 0;tag_address_2[24] <= 0;cache_block_2[24] <= 0;lru_counter_2[24] <= 0;valid_bit_3[24]  <=   0;dirty_bit_3[24] <= 0;tag_address_3[24] <= 0;cache_block_3[24] <= 0;lru_counter_3[24] <= 0;valid_bit_4[24]  <=   0;dirty_bit_4[24] <= 0;tag_address_4[24] <= 0;cache_block_4[24] <= 0;lru_counter_4[24] <= 0;
        valid_bit_1[25]  <=   0;dirty_bit_1[25] <= 0;tag_address_1[25] <= 0;cache_block_1[25] <= 0;lru_counter_1[25] <= 0;valid_bit_2[25]  <=   0;dirty_bit_2[25] <= 0;tag_address_2[25] <= 0;cache_block_2[25] <= 0;lru_counter_2[25] <= 0;valid_bit_3[25]  <=   0;dirty_bit_3[25] <= 0;tag_address_3[25] <= 0;cache_block_3[25] <= 0;lru_counter_3[25] <= 0;valid_bit_4[25]  <=   0;dirty_bit_4[25] <= 0;tag_address_4[25] <= 0;cache_block_4[25] <= 0;lru_counter_4[25] <= 0;
        valid_bit_1[26]  <=   0;dirty_bit_1[26] <= 0;tag_address_1[26] <= 0;cache_block_1[26] <= 0;lru_counter_1[26] <= 0;valid_bit_2[26]  <=   0;dirty_bit_2[26] <= 0;tag_address_2[26] <= 0;cache_block_2[26] <= 0;lru_counter_2[26] <= 0;valid_bit_3[26]  <=   0;dirty_bit_3[26] <= 0;tag_address_3[26] <= 0;cache_block_3[26] <= 0;lru_counter_3[26] <= 0;valid_bit_4[26]  <=   0;dirty_bit_4[26] <= 0;tag_address_4[26] <= 0;cache_block_4[26] <= 0;lru_counter_4[26] <= 0;
        valid_bit_1[27]  <=   0;dirty_bit_1[27] <= 0;tag_address_1[27] <= 0;cache_block_1[27] <= 0;lru_counter_1[27] <= 0;valid_bit_2[27]  <=   0;dirty_bit_2[27] <= 0;tag_address_2[27] <= 0;cache_block_2[27] <= 0;lru_counter_2[27] <= 0;valid_bit_3[27]  <=   0;dirty_bit_3[27] <= 0;tag_address_3[27] <= 0;cache_block_3[27] <= 0;lru_counter_3[27] <= 0;valid_bit_4[27]  <=   0;dirty_bit_4[27] <= 0;tag_address_4[27] <= 0;cache_block_4[27] <= 0;lru_counter_4[27] <= 0;
        valid_bit_1[28]  <=   0;dirty_bit_1[28] <= 0;tag_address_1[28] <= 0;cache_block_1[28] <= 0;lru_counter_1[28] <= 0;valid_bit_2[28]  <=   0;dirty_bit_2[28] <= 0;tag_address_2[28] <= 0;cache_block_2[28] <= 0;lru_counter_2[28] <= 0;valid_bit_3[28]  <=   0;dirty_bit_3[28] <= 0;tag_address_3[28] <= 0;cache_block_3[28] <= 0;lru_counter_3[28] <= 0;valid_bit_4[28]  <=   0;dirty_bit_4[28] <= 0;tag_address_4[28] <= 0;cache_block_4[28] <= 0;lru_counter_4[28] <= 0;
        valid_bit_1[29]  <=   0;dirty_bit_1[29] <= 0;tag_address_1[29] <= 0;cache_block_1[29] <= 0;lru_counter_1[29] <= 0;valid_bit_2[29]  <=   0;dirty_bit_2[29] <= 0;tag_address_2[29] <= 0;cache_block_2[29] <= 0;lru_counter_2[29] <= 0;valid_bit_3[29]  <=   0;dirty_bit_3[29] <= 0;tag_address_3[29] <= 0;cache_block_3[29] <= 0;lru_counter_3[29] <= 0;valid_bit_4[29]  <=   0;dirty_bit_4[29] <= 0;tag_address_4[29] <= 0;cache_block_4[29] <= 0;lru_counter_4[29] <= 0;
        valid_bit_1[30]  <=   0;dirty_bit_1[30] <= 0;tag_address_1[30] <= 0;cache_block_1[30] <= 0;lru_counter_1[30] <= 0;valid_bit_2[30]  <=   0;dirty_bit_2[30] <= 0;tag_address_2[30] <= 0;cache_block_2[30] <= 0;lru_counter_2[30] <= 0;valid_bit_3[30]  <=   0;dirty_bit_3[30] <= 0;tag_address_3[30] <= 0;cache_block_3[30] <= 0;lru_counter_3[30] <= 0;valid_bit_4[30]  <=   0;dirty_bit_4[30] <= 0;tag_address_4[30] <= 0;cache_block_4[30] <= 0;lru_counter_4[30] <= 0;
        valid_bit_1[31]  <=   0;dirty_bit_1[31] <= 0;tag_address_1[31] <= 0;cache_block_1[31] <= 0;lru_counter_1[31] <= 0;valid_bit_2[31]  <=   0;dirty_bit_2[31] <= 0;tag_address_2[31] <= 0;cache_block_2[31] <= 0;lru_counter_2[31] <= 0;valid_bit_3[31]  <=   0;dirty_bit_3[31] <= 0;tag_address_3[31] <= 0;cache_block_3[31] <= 0;lru_counter_3[31] <= 0;valid_bit_4[31]  <=   0;dirty_bit_4[31] <= 0;tag_address_4[31] <= 0;cache_block_4[31] <= 0;lru_counter_4[31] <= 0;
        valid_bit_1[32]  <=   0;dirty_bit_1[32] <= 0;tag_address_1[32] <= 0;cache_block_1[32] <= 0;lru_counter_1[32] <= 0;valid_bit_2[32]  <=   0;dirty_bit_2[32] <= 0;tag_address_2[32] <= 0;cache_block_2[32] <= 0;lru_counter_2[32] <= 0;valid_bit_3[32]  <=   0;dirty_bit_3[32] <= 0;tag_address_3[32] <= 0;cache_block_3[32] <= 0;lru_counter_3[32] <= 0;valid_bit_4[32]  <=   0;dirty_bit_4[32] <= 0;tag_address_4[32] <= 0;cache_block_4[32] <= 0;lru_counter_4[32] <= 0;
        valid_bit_1[33]  <=   0;dirty_bit_1[33] <= 0;tag_address_1[33] <= 0;cache_block_1[33] <= 0;lru_counter_1[33] <= 0;valid_bit_2[33]  <=   0;dirty_bit_2[33] <= 0;tag_address_2[33] <= 0;cache_block_2[33] <= 0;lru_counter_2[33] <= 0;valid_bit_3[33]  <=   0;dirty_bit_3[33] <= 0;tag_address_3[33] <= 0;cache_block_3[33] <= 0;lru_counter_3[33] <= 0;valid_bit_4[33]  <=   0;dirty_bit_4[33] <= 0;tag_address_4[33] <= 0;cache_block_4[33] <= 0;lru_counter_4[33] <= 0;
        valid_bit_1[34]  <=   0;dirty_bit_1[34] <= 0;tag_address_1[34] <= 0;cache_block_1[34] <= 0;lru_counter_1[34] <= 0;valid_bit_2[34]  <=   0;dirty_bit_2[34] <= 0;tag_address_2[34] <= 0;cache_block_2[34] <= 0;lru_counter_2[34] <= 0;valid_bit_3[34]  <=   0;dirty_bit_3[34] <= 0;tag_address_3[34] <= 0;cache_block_3[34] <= 0;lru_counter_3[34] <= 0;valid_bit_4[34]  <=   0;dirty_bit_4[34] <= 0;tag_address_4[34] <= 0;cache_block_4[34] <= 0;lru_counter_4[34] <= 0;
        valid_bit_1[35]  <=   0;dirty_bit_1[35] <= 0;tag_address_1[35] <= 0;cache_block_1[35] <= 0;lru_counter_1[35] <= 0;valid_bit_2[35]  <=   0;dirty_bit_2[35] <= 0;tag_address_2[35] <= 0;cache_block_2[35] <= 0;lru_counter_2[35] <= 0;valid_bit_3[35]  <=   0;dirty_bit_3[35] <= 0;tag_address_3[35] <= 0;cache_block_3[35] <= 0;lru_counter_3[35] <= 0;valid_bit_4[35]  <=   0;dirty_bit_4[35] <= 0;tag_address_4[35] <= 0;cache_block_4[35] <= 0;lru_counter_4[35] <= 0;
        valid_bit_1[36]  <=   0;dirty_bit_1[36] <= 0;tag_address_1[36] <= 0;cache_block_1[36] <= 0;lru_counter_1[36] <= 0;valid_bit_2[36]  <=   0;dirty_bit_2[36] <= 0;tag_address_2[36] <= 0;cache_block_2[36] <= 0;lru_counter_2[36] <= 0;valid_bit_3[36]  <=   0;dirty_bit_3[36] <= 0;tag_address_3[36] <= 0;cache_block_3[36] <= 0;lru_counter_3[36] <= 0;valid_bit_4[36]  <=   0;dirty_bit_4[36] <= 0;tag_address_4[36] <= 0;cache_block_4[36] <= 0;lru_counter_4[36] <= 0;
        valid_bit_1[37]  <=   0;dirty_bit_1[37] <= 0;tag_address_1[37] <= 0;cache_block_1[37] <= 0;lru_counter_1[37] <= 0;valid_bit_2[37]  <=   0;dirty_bit_2[37] <= 0;tag_address_2[37] <= 0;cache_block_2[37] <= 0;lru_counter_2[37] <= 0;valid_bit_3[37]  <=   0;dirty_bit_3[37] <= 0;tag_address_3[37] <= 0;cache_block_3[37] <= 0;lru_counter_3[37] <= 0;valid_bit_4[37]  <=   0;dirty_bit_4[37] <= 0;tag_address_4[37] <= 0;cache_block_4[37] <= 0;lru_counter_4[37] <= 0;
        valid_bit_1[38]  <=   0;dirty_bit_1[38] <= 0;tag_address_1[38] <= 0;cache_block_1[38] <= 0;lru_counter_1[38] <= 0;valid_bit_2[38]  <=   0;dirty_bit_2[38] <= 0;tag_address_2[38] <= 0;cache_block_2[38] <= 0;lru_counter_2[38] <= 0;valid_bit_3[38]  <=   0;dirty_bit_3[38] <= 0;tag_address_3[38] <= 0;cache_block_3[38] <= 0;lru_counter_3[38] <= 0;valid_bit_4[38]  <=   0;dirty_bit_4[38] <= 0;tag_address_4[38] <= 0;cache_block_4[38] <= 0;lru_counter_4[38] <= 0;
        valid_bit_1[39]  <=   0;dirty_bit_1[39] <= 0;tag_address_1[39] <= 0;cache_block_1[39] <= 0;lru_counter_1[39] <= 0;valid_bit_2[39]  <=   0;dirty_bit_2[39] <= 0;tag_address_2[39] <= 0;cache_block_2[39] <= 0;lru_counter_2[39] <= 0;valid_bit_3[39]  <=   0;dirty_bit_3[39] <= 0;tag_address_3[39] <= 0;cache_block_3[39] <= 0;lru_counter_3[39] <= 0;valid_bit_4[39]  <=   0;dirty_bit_4[39] <= 0;tag_address_4[39] <= 0;cache_block_4[39] <= 0;lru_counter_4[39] <= 0;
        valid_bit_1[40]  <=   0;dirty_bit_1[40] <= 0;tag_address_1[40] <= 0;cache_block_1[40] <= 0;lru_counter_1[40] <= 0;valid_bit_2[40]  <=   0;dirty_bit_2[40] <= 0;tag_address_2[40] <= 0;cache_block_2[40] <= 0;lru_counter_2[40] <= 0;valid_bit_3[40]  <=   0;dirty_bit_3[40] <= 0;tag_address_3[40] <= 0;cache_block_3[40] <= 0;lru_counter_3[40] <= 0;valid_bit_4[40]  <=   0;dirty_bit_4[40] <= 0;tag_address_4[40] <= 0;cache_block_4[40] <= 0;lru_counter_4[40] <= 0;
        valid_bit_1[41]  <=   0;dirty_bit_1[41] <= 0;tag_address_1[41] <= 0;cache_block_1[41] <= 0;lru_counter_1[41] <= 0;valid_bit_2[41]  <=   0;dirty_bit_2[41] <= 0;tag_address_2[41] <= 0;cache_block_2[41] <= 0;lru_counter_2[41] <= 0;valid_bit_3[41]  <=   0;dirty_bit_3[41] <= 0;tag_address_3[41] <= 0;cache_block_3[41] <= 0;lru_counter_3[41] <= 0;valid_bit_4[41]  <=   0;dirty_bit_4[41] <= 0;tag_address_4[41] <= 0;cache_block_4[41] <= 0;lru_counter_4[41] <= 0;
        valid_bit_1[42]  <=   0;dirty_bit_1[42] <= 0;tag_address_1[42] <= 0;cache_block_1[42] <= 0;lru_counter_1[42] <= 0;valid_bit_2[42]  <=   0;dirty_bit_2[42] <= 0;tag_address_2[42] <= 0;cache_block_2[42] <= 0;lru_counter_2[42] <= 0;valid_bit_3[42]  <=   0;dirty_bit_3[42] <= 0;tag_address_3[42] <= 0;cache_block_3[42] <= 0;lru_counter_3[42] <= 0;valid_bit_4[42]  <=   0;dirty_bit_4[42] <= 0;tag_address_4[42] <= 0;cache_block_4[42] <= 0;lru_counter_4[42] <= 0;
        valid_bit_1[43]  <=   0;dirty_bit_1[43] <= 0;tag_address_1[43] <= 0;cache_block_1[43] <= 0;lru_counter_1[43] <= 0;valid_bit_2[43]  <=   0;dirty_bit_2[43] <= 0;tag_address_2[43] <= 0;cache_block_2[43] <= 0;lru_counter_2[43] <= 0;valid_bit_3[43]  <=   0;dirty_bit_3[43] <= 0;tag_address_3[43] <= 0;cache_block_3[43] <= 0;lru_counter_3[43] <= 0;valid_bit_4[43]  <=   0;dirty_bit_4[43] <= 0;tag_address_4[43] <= 0;cache_block_4[43] <= 0;lru_counter_4[43] <= 0;
        valid_bit_1[44]  <=   0;dirty_bit_1[44] <= 0;tag_address_1[44] <= 0;cache_block_1[44] <= 0;lru_counter_1[44] <= 0;valid_bit_2[44]  <=   0;dirty_bit_2[44] <= 0;tag_address_2[44] <= 0;cache_block_2[44] <= 0;lru_counter_2[44] <= 0;valid_bit_3[44]  <=   0;dirty_bit_3[44] <= 0;tag_address_3[44] <= 0;cache_block_3[44] <= 0;lru_counter_3[44] <= 0;valid_bit_4[44]  <=   0;dirty_bit_4[44] <= 0;tag_address_4[44] <= 0;cache_block_4[44] <= 0;lru_counter_4[44] <= 0;
        valid_bit_1[45]  <=   0;dirty_bit_1[45] <= 0;tag_address_1[45] <= 0;cache_block_1[45] <= 0;lru_counter_1[45] <= 0;valid_bit_2[45]  <=   0;dirty_bit_2[45] <= 0;tag_address_2[45] <= 0;cache_block_2[45] <= 0;lru_counter_2[45] <= 0;valid_bit_3[45]  <=   0;dirty_bit_3[45] <= 0;tag_address_3[45] <= 0;cache_block_3[45] <= 0;lru_counter_3[45] <= 0;valid_bit_4[45]  <=   0;dirty_bit_4[45] <= 0;tag_address_4[45] <= 0;cache_block_4[45] <= 0;lru_counter_4[45] <= 0;
        valid_bit_1[46]  <=   0;dirty_bit_1[46] <= 0;tag_address_1[46] <= 0;cache_block_1[46] <= 0;lru_counter_1[46] <= 0;valid_bit_2[46]  <=   0;dirty_bit_2[46] <= 0;tag_address_2[46] <= 0;cache_block_2[46] <= 0;lru_counter_2[46] <= 0;valid_bit_3[46]  <=   0;dirty_bit_3[46] <= 0;tag_address_3[46] <= 0;cache_block_3[46] <= 0;lru_counter_3[46] <= 0;valid_bit_4[46]  <=   0;dirty_bit_4[46] <= 0;tag_address_4[46] <= 0;cache_block_4[46] <= 0;lru_counter_4[46] <= 0;
        valid_bit_1[47]  <=   0;dirty_bit_1[47] <= 0;tag_address_1[47] <= 0;cache_block_1[47] <= 0;lru_counter_1[47] <= 0;valid_bit_2[47]  <=   0;dirty_bit_2[47] <= 0;tag_address_2[47] <= 0;cache_block_2[47] <= 0;lru_counter_2[47] <= 0;valid_bit_3[47]  <=   0;dirty_bit_3[47] <= 0;tag_address_3[47] <= 0;cache_block_3[47] <= 0;lru_counter_3[47] <= 0;valid_bit_4[47]  <=   0;dirty_bit_4[47] <= 0;tag_address_4[47] <= 0;cache_block_4[47] <= 0;lru_counter_4[47] <= 0;
        valid_bit_1[48]  <=   0;dirty_bit_1[48] <= 0;tag_address_1[48] <= 0;cache_block_1[48] <= 0;lru_counter_1[48] <= 0;valid_bit_2[48]  <=   0;dirty_bit_2[48] <= 0;tag_address_2[48] <= 0;cache_block_2[48] <= 0;lru_counter_2[48] <= 0;valid_bit_3[48]  <=   0;dirty_bit_3[48] <= 0;tag_address_3[48] <= 0;cache_block_3[48] <= 0;lru_counter_3[48] <= 0;valid_bit_4[48]  <=   0;dirty_bit_4[48] <= 0;tag_address_4[48] <= 0;cache_block_4[48] <= 0;lru_counter_4[48] <= 0;
        valid_bit_1[49]  <=   0;dirty_bit_1[49] <= 0;tag_address_1[49] <= 0;cache_block_1[49] <= 0;lru_counter_1[49] <= 0;valid_bit_2[49]  <=   0;dirty_bit_2[49] <= 0;tag_address_2[49] <= 0;cache_block_2[49] <= 0;lru_counter_2[49] <= 0;valid_bit_3[49]  <=   0;dirty_bit_3[49] <= 0;tag_address_3[49] <= 0;cache_block_3[49] <= 0;lru_counter_3[49] <= 0;valid_bit_4[49]  <=   0;dirty_bit_4[49] <= 0;tag_address_4[49] <= 0;cache_block_4[49] <= 0;lru_counter_4[49] <= 0;
        valid_bit_1[50]  <=   0;dirty_bit_1[50] <= 0;tag_address_1[50] <= 0;cache_block_1[50] <= 0;lru_counter_1[50] <= 0;valid_bit_2[50]  <=   0;dirty_bit_2[50] <= 0;tag_address_2[50] <= 0;cache_block_2[50] <= 0;lru_counter_2[50] <= 0;valid_bit_3[50]  <=   0;dirty_bit_3[50] <= 0;tag_address_3[50] <= 0;cache_block_3[50] <= 0;lru_counter_3[50] <= 0;valid_bit_4[50]  <=   0;dirty_bit_4[50] <= 0;tag_address_4[50] <= 0;cache_block_4[50] <= 0;lru_counter_4[50] <= 0;
        valid_bit_1[51]  <=   0;dirty_bit_1[51] <= 0;tag_address_1[51] <= 0;cache_block_1[51] <= 0;lru_counter_1[51] <= 0;valid_bit_2[51]  <=   0;dirty_bit_2[51] <= 0;tag_address_2[51] <= 0;cache_block_2[51] <= 0;lru_counter_2[51] <= 0;valid_bit_3[51]  <=   0;dirty_bit_3[51] <= 0;tag_address_3[51] <= 0;cache_block_3[51] <= 0;lru_counter_3[51] <= 0;valid_bit_4[51]  <=   0;dirty_bit_4[51] <= 0;tag_address_4[51] <= 0;cache_block_4[51] <= 0;lru_counter_4[51] <= 0;
        valid_bit_1[52]  <=   0;dirty_bit_1[52] <= 0;tag_address_1[52] <= 0;cache_block_1[52] <= 0;lru_counter_1[52] <= 0;valid_bit_2[52]  <=   0;dirty_bit_2[52] <= 0;tag_address_2[52] <= 0;cache_block_2[52] <= 0;lru_counter_2[52] <= 0;valid_bit_3[52]  <=   0;dirty_bit_3[52] <= 0;tag_address_3[52] <= 0;cache_block_3[52] <= 0;lru_counter_3[52] <= 0;valid_bit_4[52]  <=   0;dirty_bit_4[52] <= 0;tag_address_4[52] <= 0;cache_block_4[52] <= 0;lru_counter_4[52] <= 0;
        valid_bit_1[53]  <=   0;dirty_bit_1[53] <= 0;tag_address_1[53] <= 0;cache_block_1[53] <= 0;lru_counter_1[53] <= 0;valid_bit_2[53]  <=   0;dirty_bit_2[53] <= 0;tag_address_2[53] <= 0;cache_block_2[53] <= 0;lru_counter_2[53] <= 0;valid_bit_3[53]  <=   0;dirty_bit_3[53] <= 0;tag_address_3[53] <= 0;cache_block_3[53] <= 0;lru_counter_3[53] <= 0;valid_bit_4[53]  <=   0;dirty_bit_4[53] <= 0;tag_address_4[53] <= 0;cache_block_4[53] <= 0;lru_counter_4[53] <= 0;
        valid_bit_1[54]  <=   0;dirty_bit_1[54] <= 0;tag_address_1[54] <= 0;cache_block_1[54] <= 0;lru_counter_1[54] <= 0;valid_bit_2[54]  <=   0;dirty_bit_2[54] <= 0;tag_address_2[54] <= 0;cache_block_2[54] <= 0;lru_counter_2[54] <= 0;valid_bit_3[54]  <=   0;dirty_bit_3[54] <= 0;tag_address_3[54] <= 0;cache_block_3[54] <= 0;lru_counter_3[54] <= 0;valid_bit_4[54]  <=   0;dirty_bit_4[54] <= 0;tag_address_4[54] <= 0;cache_block_4[54] <= 0;lru_counter_4[54] <= 0;
        valid_bit_1[55]  <=   0;dirty_bit_1[55] <= 0;tag_address_1[55] <= 0;cache_block_1[55] <= 0;lru_counter_1[55] <= 0;valid_bit_2[55]  <=   0;dirty_bit_2[55] <= 0;tag_address_2[55] <= 0;cache_block_2[55] <= 0;lru_counter_2[55] <= 0;valid_bit_3[55]  <=   0;dirty_bit_3[55] <= 0;tag_address_3[55] <= 0;cache_block_3[55] <= 0;lru_counter_3[55] <= 0;valid_bit_4[55]  <=   0;dirty_bit_4[55] <= 0;tag_address_4[55] <= 0;cache_block_4[55] <= 0;lru_counter_4[55] <= 0;
        valid_bit_1[56]  <=   0;dirty_bit_1[56] <= 0;tag_address_1[56] <= 0;cache_block_1[56] <= 0;lru_counter_1[56] <= 0;valid_bit_2[56]  <=   0;dirty_bit_2[56] <= 0;tag_address_2[56] <= 0;cache_block_2[56] <= 0;lru_counter_2[56] <= 0;valid_bit_3[56]  <=   0;dirty_bit_3[56] <= 0;tag_address_3[56] <= 0;cache_block_3[56] <= 0;lru_counter_3[56] <= 0;valid_bit_4[56]  <=   0;dirty_bit_4[56] <= 0;tag_address_4[56] <= 0;cache_block_4[56] <= 0;lru_counter_4[56] <= 0;
        valid_bit_1[57]  <=   0;dirty_bit_1[57] <= 0;tag_address_1[57] <= 0;cache_block_1[57] <= 0;lru_counter_1[57] <= 0;valid_bit_2[57]  <=   0;dirty_bit_2[57] <= 0;tag_address_2[57] <= 0;cache_block_2[57] <= 0;lru_counter_2[57] <= 0;valid_bit_3[57]  <=   0;dirty_bit_3[57] <= 0;tag_address_3[57] <= 0;cache_block_3[57] <= 0;lru_counter_3[57] <= 0;valid_bit_4[57]  <=   0;dirty_bit_4[57] <= 0;tag_address_4[57] <= 0;cache_block_4[57] <= 0;lru_counter_4[57] <= 0;
        valid_bit_1[58]  <=   0;dirty_bit_1[58] <= 0;tag_address_1[58] <= 0;cache_block_1[58] <= 0;lru_counter_1[58] <= 0;valid_bit_2[58]  <=   0;dirty_bit_2[58] <= 0;tag_address_2[58] <= 0;cache_block_2[58] <= 0;lru_counter_2[58] <= 0;valid_bit_3[58]  <=   0;dirty_bit_3[58] <= 0;tag_address_3[58] <= 0;cache_block_3[58] <= 0;lru_counter_3[58] <= 0;valid_bit_4[58]  <=   0;dirty_bit_4[58] <= 0;tag_address_4[58] <= 0;cache_block_4[58] <= 0;lru_counter_4[58] <= 0;
        valid_bit_1[59]  <=   0;dirty_bit_1[59] <= 0;tag_address_1[59] <= 0;cache_block_1[59] <= 0;lru_counter_1[59] <= 0;valid_bit_2[59]  <=   0;dirty_bit_2[59] <= 0;tag_address_2[59] <= 0;cache_block_2[59] <= 0;lru_counter_2[59] <= 0;valid_bit_3[59]  <=   0;dirty_bit_3[59] <= 0;tag_address_3[59] <= 0;cache_block_3[59] <= 0;lru_counter_3[59] <= 0;valid_bit_4[59]  <=   0;dirty_bit_4[59] <= 0;tag_address_4[59] <= 0;cache_block_4[59] <= 0;lru_counter_4[59] <= 0;
        valid_bit_1[60]  <=   0;dirty_bit_1[60] <= 0;tag_address_1[60] <= 0;cache_block_1[60] <= 0;lru_counter_1[60] <= 0;valid_bit_2[60]  <=   0;dirty_bit_2[60] <= 0;tag_address_2[60] <= 0;cache_block_2[60] <= 0;lru_counter_2[60] <= 0;valid_bit_3[60]  <=   0;dirty_bit_3[60] <= 0;tag_address_3[60] <= 0;cache_block_3[60] <= 0;lru_counter_3[60] <= 0;valid_bit_4[60]  <=   0;dirty_bit_4[60] <= 0;tag_address_4[60] <= 0;cache_block_4[60] <= 0;lru_counter_4[60] <= 0;
        valid_bit_1[61]  <=   0;dirty_bit_1[61] <= 0;tag_address_1[61] <= 0;cache_block_1[61] <= 0;lru_counter_1[61] <= 0;valid_bit_2[61]  <=   0;dirty_bit_2[61] <= 0;tag_address_2[61] <= 0;cache_block_2[61] <= 0;lru_counter_2[61] <= 0;valid_bit_3[61]  <=   0;dirty_bit_3[61] <= 0;tag_address_3[61] <= 0;cache_block_3[61] <= 0;lru_counter_3[61] <= 0;valid_bit_4[61]  <=   0;dirty_bit_4[61] <= 0;tag_address_4[61] <= 0;cache_block_4[61] <= 0;lru_counter_4[61] <= 0;
        valid_bit_1[62]  <=   0;dirty_bit_1[62] <= 0;tag_address_1[62] <= 0;cache_block_1[62] <= 0;lru_counter_1[62] <= 0;valid_bit_2[62]  <=   0;dirty_bit_2[62] <= 0;tag_address_2[62] <= 0;cache_block_2[62] <= 0;lru_counter_2[62] <= 0;valid_bit_3[62]  <=   0;dirty_bit_3[62] <= 0;tag_address_3[62] <= 0;cache_block_3[62] <= 0;lru_counter_3[62] <= 0;valid_bit_4[62]  <=   0;dirty_bit_4[62] <= 0;tag_address_4[62] <= 0;cache_block_4[62] <= 0;lru_counter_4[62] <= 0;
        valid_bit_1[63]  <=   0;dirty_bit_1[63] <= 0;tag_address_1[63] <= 0;cache_block_1[63] <= 0;lru_counter_1[63] <= 0;valid_bit_2[63]  <=   0;dirty_bit_2[63] <= 0;tag_address_2[63] <= 0;cache_block_2[63] <= 0;lru_counter_2[63] <= 0;valid_bit_3[63]  <=   0;dirty_bit_3[63] <= 0;tag_address_3[63] <= 0;cache_block_3[63] <= 0;lru_counter_3[63] <= 0;valid_bit_4[63]  <=   0;dirty_bit_4[63] <= 0;tag_address_4[63] <= 0;cache_block_4[63] <= 0;lru_counter_4[63] <= 0;
        valid_bit_1[64]  <=   0;dirty_bit_1[64] <= 0;tag_address_1[64] <= 0;cache_block_1[64] <= 0;lru_counter_1[64] <= 0;valid_bit_2[64]  <=   0;dirty_bit_2[64] <= 0;tag_address_2[64] <= 0;cache_block_2[64] <= 0;lru_counter_2[64] <= 0;valid_bit_3[64]  <=   0;dirty_bit_3[64] <= 0;tag_address_3[64] <= 0;cache_block_3[64] <= 0;lru_counter_3[64] <= 0;valid_bit_4[64]  <=   0;dirty_bit_4[64] <= 0;tag_address_4[64] <= 0;cache_block_4[64] <= 0;lru_counter_4[64] <= 0;
        valid_bit_1[65]  <=   0;dirty_bit_1[65] <= 0;tag_address_1[65] <= 0;cache_block_1[65] <= 0;lru_counter_1[65] <= 0;valid_bit_2[65]  <=   0;dirty_bit_2[65] <= 0;tag_address_2[65] <= 0;cache_block_2[65] <= 0;lru_counter_2[65] <= 0;valid_bit_3[65]  <=   0;dirty_bit_3[65] <= 0;tag_address_3[65] <= 0;cache_block_3[65] <= 0;lru_counter_3[65] <= 0;valid_bit_4[65]  <=   0;dirty_bit_4[65] <= 0;tag_address_4[65] <= 0;cache_block_4[65] <= 0;lru_counter_4[65] <= 0;
        valid_bit_1[66]  <=   0;dirty_bit_1[66] <= 0;tag_address_1[66] <= 0;cache_block_1[66] <= 0;lru_counter_1[66] <= 0;valid_bit_2[66]  <=   0;dirty_bit_2[66] <= 0;tag_address_2[66] <= 0;cache_block_2[66] <= 0;lru_counter_2[66] <= 0;valid_bit_3[66]  <=   0;dirty_bit_3[66] <= 0;tag_address_3[66] <= 0;cache_block_3[66] <= 0;lru_counter_3[66] <= 0;valid_bit_4[66]  <=   0;dirty_bit_4[66] <= 0;tag_address_4[66] <= 0;cache_block_4[66] <= 0;lru_counter_4[66] <= 0;
        valid_bit_1[67]  <=   0;dirty_bit_1[67] <= 0;tag_address_1[67] <= 0;cache_block_1[67] <= 0;lru_counter_1[67] <= 0;valid_bit_2[67]  <=   0;dirty_bit_2[67] <= 0;tag_address_2[67] <= 0;cache_block_2[67] <= 0;lru_counter_2[67] <= 0;valid_bit_3[67]  <=   0;dirty_bit_3[67] <= 0;tag_address_3[67] <= 0;cache_block_3[67] <= 0;lru_counter_3[67] <= 0;valid_bit_4[67]  <=   0;dirty_bit_4[67] <= 0;tag_address_4[67] <= 0;cache_block_4[67] <= 0;lru_counter_4[67] <= 0;
        valid_bit_1[68]  <=   0;dirty_bit_1[68] <= 0;tag_address_1[68] <= 0;cache_block_1[68] <= 0;lru_counter_1[68] <= 0;valid_bit_2[68]  <=   0;dirty_bit_2[68] <= 0;tag_address_2[68] <= 0;cache_block_2[68] <= 0;lru_counter_2[68] <= 0;valid_bit_3[68]  <=   0;dirty_bit_3[68] <= 0;tag_address_3[68] <= 0;cache_block_3[68] <= 0;lru_counter_3[68] <= 0;valid_bit_4[68]  <=   0;dirty_bit_4[68] <= 0;tag_address_4[68] <= 0;cache_block_4[68] <= 0;lru_counter_4[68] <= 0;
        valid_bit_1[69]  <=   0;dirty_bit_1[69] <= 0;tag_address_1[69] <= 0;cache_block_1[69] <= 0;lru_counter_1[69] <= 0;valid_bit_2[69]  <=   0;dirty_bit_2[69] <= 0;tag_address_2[69] <= 0;cache_block_2[69] <= 0;lru_counter_2[69] <= 0;valid_bit_3[69]  <=   0;dirty_bit_3[69] <= 0;tag_address_3[69] <= 0;cache_block_3[69] <= 0;lru_counter_3[69] <= 0;valid_bit_4[69]  <=   0;dirty_bit_4[69] <= 0;tag_address_4[69] <= 0;cache_block_4[69] <= 0;lru_counter_4[69] <= 0;
        valid_bit_1[70]  <=   0;dirty_bit_1[70] <= 0;tag_address_1[70] <= 0;cache_block_1[70] <= 0;lru_counter_1[70] <= 0;valid_bit_2[70]  <=   0;dirty_bit_2[70] <= 0;tag_address_2[70] <= 0;cache_block_2[70] <= 0;lru_counter_2[70] <= 0;valid_bit_3[70]  <=   0;dirty_bit_3[70] <= 0;tag_address_3[70] <= 0;cache_block_3[70] <= 0;lru_counter_3[70] <= 0;valid_bit_4[70]  <=   0;dirty_bit_4[70] <= 0;tag_address_4[70] <= 0;cache_block_4[70] <= 0;lru_counter_4[70] <= 0;
        valid_bit_1[71]  <=   0;dirty_bit_1[71] <= 0;tag_address_1[71] <= 0;cache_block_1[71] <= 0;lru_counter_1[71] <= 0;valid_bit_2[71]  <=   0;dirty_bit_2[71] <= 0;tag_address_2[71] <= 0;cache_block_2[71] <= 0;lru_counter_2[71] <= 0;valid_bit_3[71]  <=   0;dirty_bit_3[71] <= 0;tag_address_3[71] <= 0;cache_block_3[71] <= 0;lru_counter_3[71] <= 0;valid_bit_4[71]  <=   0;dirty_bit_4[71] <= 0;tag_address_4[71] <= 0;cache_block_4[71] <= 0;lru_counter_4[71] <= 0;
        valid_bit_1[72]  <=   0;dirty_bit_1[72] <= 0;tag_address_1[72] <= 0;cache_block_1[72] <= 0;lru_counter_1[72] <= 0;valid_bit_2[72]  <=   0;dirty_bit_2[72] <= 0;tag_address_2[72] <= 0;cache_block_2[72] <= 0;lru_counter_2[72] <= 0;valid_bit_3[72]  <=   0;dirty_bit_3[72] <= 0;tag_address_3[72] <= 0;cache_block_3[72] <= 0;lru_counter_3[72] <= 0;valid_bit_4[72]  <=   0;dirty_bit_4[72] <= 0;tag_address_4[72] <= 0;cache_block_4[72] <= 0;lru_counter_4[72] <= 0;
        valid_bit_1[73]  <=   0;dirty_bit_1[73] <= 0;tag_address_1[73] <= 0;cache_block_1[73] <= 0;lru_counter_1[73] <= 0;valid_bit_2[73]  <=   0;dirty_bit_2[73] <= 0;tag_address_2[73] <= 0;cache_block_2[73] <= 0;lru_counter_2[73] <= 0;valid_bit_3[73]  <=   0;dirty_bit_3[73] <= 0;tag_address_3[73] <= 0;cache_block_3[73] <= 0;lru_counter_3[73] <= 0;valid_bit_4[73]  <=   0;dirty_bit_4[73] <= 0;tag_address_4[73] <= 0;cache_block_4[73] <= 0;lru_counter_4[73] <= 0;
        valid_bit_1[74]  <=   0;dirty_bit_1[74] <= 0;tag_address_1[74] <= 0;cache_block_1[74] <= 0;lru_counter_1[74] <= 0;valid_bit_2[74]  <=   0;dirty_bit_2[74] <= 0;tag_address_2[74] <= 0;cache_block_2[74] <= 0;lru_counter_2[74] <= 0;valid_bit_3[74]  <=   0;dirty_bit_3[74] <= 0;tag_address_3[74] <= 0;cache_block_3[74] <= 0;lru_counter_3[74] <= 0;valid_bit_4[74]  <=   0;dirty_bit_4[74] <= 0;tag_address_4[74] <= 0;cache_block_4[74] <= 0;lru_counter_4[74] <= 0;
        valid_bit_1[75]  <=   0;dirty_bit_1[75] <= 0;tag_address_1[75] <= 0;cache_block_1[75] <= 0;lru_counter_1[75] <= 0;valid_bit_2[75]  <=   0;dirty_bit_2[75] <= 0;tag_address_2[75] <= 0;cache_block_2[75] <= 0;lru_counter_2[75] <= 0;valid_bit_3[75]  <=   0;dirty_bit_3[75] <= 0;tag_address_3[75] <= 0;cache_block_3[75] <= 0;lru_counter_3[75] <= 0;valid_bit_4[75]  <=   0;dirty_bit_4[75] <= 0;tag_address_4[75] <= 0;cache_block_4[75] <= 0;lru_counter_4[75] <= 0;
        valid_bit_1[76]  <=   0;dirty_bit_1[76] <= 0;tag_address_1[76] <= 0;cache_block_1[76] <= 0;lru_counter_1[76] <= 0;valid_bit_2[76]  <=   0;dirty_bit_2[76] <= 0;tag_address_2[76] <= 0;cache_block_2[76] <= 0;lru_counter_2[76] <= 0;valid_bit_3[76]  <=   0;dirty_bit_3[76] <= 0;tag_address_3[76] <= 0;cache_block_3[76] <= 0;lru_counter_3[76] <= 0;valid_bit_4[76]  <=   0;dirty_bit_4[76] <= 0;tag_address_4[76] <= 0;cache_block_4[76] <= 0;lru_counter_4[76] <= 0;
        valid_bit_1[77]  <=   0;dirty_bit_1[77] <= 0;tag_address_1[77] <= 0;cache_block_1[77] <= 0;lru_counter_1[77] <= 0;valid_bit_2[77]  <=   0;dirty_bit_2[77] <= 0;tag_address_2[77] <= 0;cache_block_2[77] <= 0;lru_counter_2[77] <= 0;valid_bit_3[77]  <=   0;dirty_bit_3[77] <= 0;tag_address_3[77] <= 0;cache_block_3[77] <= 0;lru_counter_3[77] <= 0;valid_bit_4[77]  <=   0;dirty_bit_4[77] <= 0;tag_address_4[77] <= 0;cache_block_4[77] <= 0;lru_counter_4[77] <= 0;
        valid_bit_1[78]  <=   0;dirty_bit_1[78] <= 0;tag_address_1[78] <= 0;cache_block_1[78] <= 0;lru_counter_1[78] <= 0;valid_bit_2[78]  <=   0;dirty_bit_2[78] <= 0;tag_address_2[78] <= 0;cache_block_2[78] <= 0;lru_counter_2[78] <= 0;valid_bit_3[78]  <=   0;dirty_bit_3[78] <= 0;tag_address_3[78] <= 0;cache_block_3[78] <= 0;lru_counter_3[78] <= 0;valid_bit_4[78]  <=   0;dirty_bit_4[78] <= 0;tag_address_4[78] <= 0;cache_block_4[78] <= 0;lru_counter_4[78] <= 0;
        valid_bit_1[79]  <=   0;dirty_bit_1[79] <= 0;tag_address_1[79] <= 0;cache_block_1[79] <= 0;lru_counter_1[79] <= 0;valid_bit_2[79]  <=   0;dirty_bit_2[79] <= 0;tag_address_2[79] <= 0;cache_block_2[79] <= 0;lru_counter_2[79] <= 0;valid_bit_3[79]  <=   0;dirty_bit_3[79] <= 0;tag_address_3[79] <= 0;cache_block_3[79] <= 0;lru_counter_3[79] <= 0;valid_bit_4[79]  <=   0;dirty_bit_4[79] <= 0;tag_address_4[79] <= 0;cache_block_4[79] <= 0;lru_counter_4[79] <= 0;
        valid_bit_1[80]  <=   0;dirty_bit_1[80] <= 0;tag_address_1[80] <= 0;cache_block_1[80] <= 0;lru_counter_1[80] <= 0;valid_bit_2[80]  <=   0;dirty_bit_2[80] <= 0;tag_address_2[80] <= 0;cache_block_2[80] <= 0;lru_counter_2[80] <= 0;valid_bit_3[80]  <=   0;dirty_bit_3[80] <= 0;tag_address_3[80] <= 0;cache_block_3[80] <= 0;lru_counter_3[80] <= 0;valid_bit_4[80]  <=   0;dirty_bit_4[80] <= 0;tag_address_4[80] <= 0;cache_block_4[80] <= 0;lru_counter_4[80] <= 0;
        valid_bit_1[81]  <=   0;dirty_bit_1[81] <= 0;tag_address_1[81] <= 0;cache_block_1[81] <= 0;lru_counter_1[81] <= 0;valid_bit_2[81]  <=   0;dirty_bit_2[81] <= 0;tag_address_2[81] <= 0;cache_block_2[81] <= 0;lru_counter_2[81] <= 0;valid_bit_3[81]  <=   0;dirty_bit_3[81] <= 0;tag_address_3[81] <= 0;cache_block_3[81] <= 0;lru_counter_3[81] <= 0;valid_bit_4[81]  <=   0;dirty_bit_4[81] <= 0;tag_address_4[81] <= 0;cache_block_4[81] <= 0;lru_counter_4[81] <= 0;
        valid_bit_1[82]  <=   0;dirty_bit_1[82] <= 0;tag_address_1[82] <= 0;cache_block_1[82] <= 0;lru_counter_1[82] <= 0;valid_bit_2[82]  <=   0;dirty_bit_2[82] <= 0;tag_address_2[82] <= 0;cache_block_2[82] <= 0;lru_counter_2[82] <= 0;valid_bit_3[82]  <=   0;dirty_bit_3[82] <= 0;tag_address_3[82] <= 0;cache_block_3[82] <= 0;lru_counter_3[82] <= 0;valid_bit_4[82]  <=   0;dirty_bit_4[82] <= 0;tag_address_4[82] <= 0;cache_block_4[82] <= 0;lru_counter_4[82] <= 0;
        valid_bit_1[83]  <=   0;dirty_bit_1[83] <= 0;tag_address_1[83] <= 0;cache_block_1[83] <= 0;lru_counter_1[83] <= 0;valid_bit_2[83]  <=   0;dirty_bit_2[83] <= 0;tag_address_2[83] <= 0;cache_block_2[83] <= 0;lru_counter_2[83] <= 0;valid_bit_3[83]  <=   0;dirty_bit_3[83] <= 0;tag_address_3[83] <= 0;cache_block_3[83] <= 0;lru_counter_3[83] <= 0;valid_bit_4[83]  <=   0;dirty_bit_4[83] <= 0;tag_address_4[83] <= 0;cache_block_4[83] <= 0;lru_counter_4[83] <= 0;
        valid_bit_1[84]  <=   0;dirty_bit_1[84] <= 0;tag_address_1[84] <= 0;cache_block_1[84] <= 0;lru_counter_1[84] <= 0;valid_bit_2[84]  <=   0;dirty_bit_2[84] <= 0;tag_address_2[84] <= 0;cache_block_2[84] <= 0;lru_counter_2[84] <= 0;valid_bit_3[84]  <=   0;dirty_bit_3[84] <= 0;tag_address_3[84] <= 0;cache_block_3[84] <= 0;lru_counter_3[84] <= 0;valid_bit_4[84]  <=   0;dirty_bit_4[84] <= 0;tag_address_4[84] <= 0;cache_block_4[84] <= 0;lru_counter_4[84] <= 0;
        valid_bit_1[85]  <=   0;dirty_bit_1[85] <= 0;tag_address_1[85] <= 0;cache_block_1[85] <= 0;lru_counter_1[85] <= 0;valid_bit_2[85]  <=   0;dirty_bit_2[85] <= 0;tag_address_2[85] <= 0;cache_block_2[85] <= 0;lru_counter_2[85] <= 0;valid_bit_3[85]  <=   0;dirty_bit_3[85] <= 0;tag_address_3[85] <= 0;cache_block_3[85] <= 0;lru_counter_3[85] <= 0;valid_bit_4[85]  <=   0;dirty_bit_4[85] <= 0;tag_address_4[85] <= 0;cache_block_4[85] <= 0;lru_counter_4[85] <= 0;
        valid_bit_1[86]  <=   0;dirty_bit_1[86] <= 0;tag_address_1[86] <= 0;cache_block_1[86] <= 0;lru_counter_1[86] <= 0;valid_bit_2[86]  <=   0;dirty_bit_2[86] <= 0;tag_address_2[86] <= 0;cache_block_2[86] <= 0;lru_counter_2[86] <= 0;valid_bit_3[86]  <=   0;dirty_bit_3[86] <= 0;tag_address_3[86] <= 0;cache_block_3[86] <= 0;lru_counter_3[86] <= 0;valid_bit_4[86]  <=   0;dirty_bit_4[86] <= 0;tag_address_4[86] <= 0;cache_block_4[86] <= 0;lru_counter_4[86] <= 0;
        valid_bit_1[87]  <=   0;dirty_bit_1[87] <= 0;tag_address_1[87] <= 0;cache_block_1[87] <= 0;lru_counter_1[87] <= 0;valid_bit_2[87]  <=   0;dirty_bit_2[87] <= 0;tag_address_2[87] <= 0;cache_block_2[87] <= 0;lru_counter_2[87] <= 0;valid_bit_3[87]  <=   0;dirty_bit_3[87] <= 0;tag_address_3[87] <= 0;cache_block_3[87] <= 0;lru_counter_3[87] <= 0;valid_bit_4[87]  <=   0;dirty_bit_4[87] <= 0;tag_address_4[87] <= 0;cache_block_4[87] <= 0;lru_counter_4[87] <= 0;
        valid_bit_1[88]  <=   0;dirty_bit_1[88] <= 0;tag_address_1[88] <= 0;cache_block_1[88] <= 0;lru_counter_1[88] <= 0;valid_bit_2[88]  <=   0;dirty_bit_2[88] <= 0;tag_address_2[88] <= 0;cache_block_2[88] <= 0;lru_counter_2[88] <= 0;valid_bit_3[88]  <=   0;dirty_bit_3[88] <= 0;tag_address_3[88] <= 0;cache_block_3[88] <= 0;lru_counter_3[88] <= 0;valid_bit_4[88]  <=   0;dirty_bit_4[88] <= 0;tag_address_4[88] <= 0;cache_block_4[88] <= 0;lru_counter_4[88] <= 0;
        valid_bit_1[89]  <=   0;dirty_bit_1[89] <= 0;tag_address_1[89] <= 0;cache_block_1[89] <= 0;lru_counter_1[89] <= 0;valid_bit_2[89]  <=   0;dirty_bit_2[89] <= 0;tag_address_2[89] <= 0;cache_block_2[89] <= 0;lru_counter_2[89] <= 0;valid_bit_3[89]  <=   0;dirty_bit_3[89] <= 0;tag_address_3[89] <= 0;cache_block_3[89] <= 0;lru_counter_3[89] <= 0;valid_bit_4[89]  <=   0;dirty_bit_4[89] <= 0;tag_address_4[89] <= 0;cache_block_4[89] <= 0;lru_counter_4[89] <= 0;
        valid_bit_1[90]  <=   0;dirty_bit_1[90] <= 0;tag_address_1[90] <= 0;cache_block_1[90] <= 0;lru_counter_1[90] <= 0;valid_bit_2[90]  <=   0;dirty_bit_2[90] <= 0;tag_address_2[90] <= 0;cache_block_2[90] <= 0;lru_counter_2[90] <= 0;valid_bit_3[90]  <=   0;dirty_bit_3[90] <= 0;tag_address_3[90] <= 0;cache_block_3[90] <= 0;lru_counter_3[90] <= 0;valid_bit_4[90]  <=   0;dirty_bit_4[90] <= 0;tag_address_4[90] <= 0;cache_block_4[90] <= 0;lru_counter_4[90] <= 0;
        valid_bit_1[91]  <=   0;dirty_bit_1[91] <= 0;tag_address_1[91] <= 0;cache_block_1[91] <= 0;lru_counter_1[91] <= 0;valid_bit_2[91]  <=   0;dirty_bit_2[91] <= 0;tag_address_2[91] <= 0;cache_block_2[91] <= 0;lru_counter_2[91] <= 0;valid_bit_3[91]  <=   0;dirty_bit_3[91] <= 0;tag_address_3[91] <= 0;cache_block_3[91] <= 0;lru_counter_3[91] <= 0;valid_bit_4[91]  <=   0;dirty_bit_4[91] <= 0;tag_address_4[91] <= 0;cache_block_4[91] <= 0;lru_counter_4[91] <= 0;
        valid_bit_1[92]  <=   0;dirty_bit_1[92] <= 0;tag_address_1[92] <= 0;cache_block_1[92] <= 0;lru_counter_1[92] <= 0;valid_bit_2[92]  <=   0;dirty_bit_2[92] <= 0;tag_address_2[92] <= 0;cache_block_2[92] <= 0;lru_counter_2[92] <= 0;valid_bit_3[92]  <=   0;dirty_bit_3[92] <= 0;tag_address_3[92] <= 0;cache_block_3[92] <= 0;lru_counter_3[92] <= 0;valid_bit_4[92]  <=   0;dirty_bit_4[92] <= 0;tag_address_4[92] <= 0;cache_block_4[92] <= 0;lru_counter_4[92] <= 0;
        valid_bit_1[93]  <=   0;dirty_bit_1[93] <= 0;tag_address_1[93] <= 0;cache_block_1[93] <= 0;lru_counter_1[93] <= 0;valid_bit_2[93]  <=   0;dirty_bit_2[93] <= 0;tag_address_2[93] <= 0;cache_block_2[93] <= 0;lru_counter_2[93] <= 0;valid_bit_3[93]  <=   0;dirty_bit_3[93] <= 0;tag_address_3[93] <= 0;cache_block_3[93] <= 0;lru_counter_3[93] <= 0;valid_bit_4[93]  <=   0;dirty_bit_4[93] <= 0;tag_address_4[93] <= 0;cache_block_4[93] <= 0;lru_counter_4[93] <= 0;
        valid_bit_1[94]  <=   0;dirty_bit_1[94] <= 0;tag_address_1[94] <= 0;cache_block_1[94] <= 0;lru_counter_1[94] <= 0;valid_bit_2[94]  <=   0;dirty_bit_2[94] <= 0;tag_address_2[94] <= 0;cache_block_2[94] <= 0;lru_counter_2[94] <= 0;valid_bit_3[94]  <=   0;dirty_bit_3[94] <= 0;tag_address_3[94] <= 0;cache_block_3[94] <= 0;lru_counter_3[94] <= 0;valid_bit_4[94]  <=   0;dirty_bit_4[94] <= 0;tag_address_4[94] <= 0;cache_block_4[94] <= 0;lru_counter_4[94] <= 0;
        valid_bit_1[95]  <=   0;dirty_bit_1[95] <= 0;tag_address_1[95] <= 0;cache_block_1[95] <= 0;lru_counter_1[95] <= 0;valid_bit_2[95]  <=   0;dirty_bit_2[95] <= 0;tag_address_2[95] <= 0;cache_block_2[95] <= 0;lru_counter_2[95] <= 0;valid_bit_3[95]  <=   0;dirty_bit_3[95] <= 0;tag_address_3[95] <= 0;cache_block_3[95] <= 0;lru_counter_3[95] <= 0;valid_bit_4[95]  <=   0;dirty_bit_4[95] <= 0;tag_address_4[95] <= 0;cache_block_4[95] <= 0;lru_counter_4[95] <= 0;
        valid_bit_1[96]  <=   0;dirty_bit_1[96] <= 0;tag_address_1[96] <= 0;cache_block_1[96] <= 0;lru_counter_1[96] <= 0;valid_bit_2[96]  <=   0;dirty_bit_2[96] <= 0;tag_address_2[96] <= 0;cache_block_2[96] <= 0;lru_counter_2[96] <= 0;valid_bit_3[96]  <=   0;dirty_bit_3[96] <= 0;tag_address_3[96] <= 0;cache_block_3[96] <= 0;lru_counter_3[96] <= 0;valid_bit_4[96]  <=   0;dirty_bit_4[96] <= 0;tag_address_4[96] <= 0;cache_block_4[96] <= 0;lru_counter_4[96] <= 0;
        valid_bit_1[97]  <=   0;dirty_bit_1[97] <= 0;tag_address_1[97] <= 0;cache_block_1[97] <= 0;lru_counter_1[97] <= 0;valid_bit_2[97]  <=   0;dirty_bit_2[97] <= 0;tag_address_2[97] <= 0;cache_block_2[97] <= 0;lru_counter_2[97] <= 0;valid_bit_3[97]  <=   0;dirty_bit_3[97] <= 0;tag_address_3[97] <= 0;cache_block_3[97] <= 0;lru_counter_3[97] <= 0;valid_bit_4[97]  <=   0;dirty_bit_4[97] <= 0;tag_address_4[97] <= 0;cache_block_4[97] <= 0;lru_counter_4[97] <= 0;
        valid_bit_1[98]  <=   0;dirty_bit_1[98] <= 0;tag_address_1[98] <= 0;cache_block_1[98] <= 0;lru_counter_1[98] <= 0;valid_bit_2[98]  <=   0;dirty_bit_2[98] <= 0;tag_address_2[98] <= 0;cache_block_2[98] <= 0;lru_counter_2[98] <= 0;valid_bit_3[98]  <=   0;dirty_bit_3[98] <= 0;tag_address_3[98] <= 0;cache_block_3[98] <= 0;lru_counter_3[98] <= 0;valid_bit_4[98]  <=   0;dirty_bit_4[98] <= 0;tag_address_4[98] <= 0;cache_block_4[98] <= 0;lru_counter_4[98] <= 0;
        valid_bit_1[99]  <=   0;dirty_bit_1[99] <= 0;tag_address_1[99] <= 0;cache_block_1[99] <= 0;lru_counter_1[99] <= 0;valid_bit_2[99]  <=   0;dirty_bit_2[99] <= 0;tag_address_2[99] <= 0;cache_block_2[99] <= 0;lru_counter_2[99] <= 0;valid_bit_3[99]  <=   0;dirty_bit_3[99] <= 0;tag_address_3[99] <= 0;cache_block_3[99] <= 0;lru_counter_3[99] <= 0;valid_bit_4[99]  <=   0;dirty_bit_4[99] <= 0;tag_address_4[99] <= 0;cache_block_4[99] <= 0;lru_counter_4[99] <= 0;
        valid_bit_1[100]  <=   0;dirty_bit_1[100] <= 0;tag_address_1[100] <= 0;cache_block_1[100] <= 0;lru_counter_1[100] <= 0;valid_bit_2[100]  <=   0;dirty_bit_2[100] <= 0;tag_address_2[100] <= 0;cache_block_2[100] <= 0;lru_counter_2[100] <= 0;valid_bit_3[100]  <=   0;dirty_bit_3[100] <= 0;tag_address_3[100] <= 0;cache_block_3[100] <= 0;lru_counter_3[100] <= 0;valid_bit_4[100]  <=   0;dirty_bit_4[100] <= 0;tag_address_4[100] <= 0;cache_block_4[100] <= 0;lru_counter_4[100] <= 0;
        valid_bit_1[101]  <=   0;dirty_bit_1[101] <= 0;tag_address_1[101] <= 0;cache_block_1[101] <= 0;lru_counter_1[101] <= 0;valid_bit_2[101]  <=   0;dirty_bit_2[101] <= 0;tag_address_2[101] <= 0;cache_block_2[101] <= 0;lru_counter_2[101] <= 0;valid_bit_3[101]  <=   0;dirty_bit_3[101] <= 0;tag_address_3[101] <= 0;cache_block_3[101] <= 0;lru_counter_3[101] <= 0;valid_bit_4[101]  <=   0;dirty_bit_4[101] <= 0;tag_address_4[101] <= 0;cache_block_4[101] <= 0;lru_counter_4[101] <= 0;
        valid_bit_1[102]  <=   0;dirty_bit_1[102] <= 0;tag_address_1[102] <= 0;cache_block_1[102] <= 0;lru_counter_1[102] <= 0;valid_bit_2[102]  <=   0;dirty_bit_2[102] <= 0;tag_address_2[102] <= 0;cache_block_2[102] <= 0;lru_counter_2[102] <= 0;valid_bit_3[102]  <=   0;dirty_bit_3[102] <= 0;tag_address_3[102] <= 0;cache_block_3[102] <= 0;lru_counter_3[102] <= 0;valid_bit_4[102]  <=   0;dirty_bit_4[102] <= 0;tag_address_4[102] <= 0;cache_block_4[102] <= 0;lru_counter_4[102] <= 0;
        valid_bit_1[103]  <=   0;dirty_bit_1[103] <= 0;tag_address_1[103] <= 0;cache_block_1[103] <= 0;lru_counter_1[103] <= 0;valid_bit_2[103]  <=   0;dirty_bit_2[103] <= 0;tag_address_2[103] <= 0;cache_block_2[103] <= 0;lru_counter_2[103] <= 0;valid_bit_3[103]  <=   0;dirty_bit_3[103] <= 0;tag_address_3[103] <= 0;cache_block_3[103] <= 0;lru_counter_3[103] <= 0;valid_bit_4[103]  <=   0;dirty_bit_4[103] <= 0;tag_address_4[103] <= 0;cache_block_4[103] <= 0;lru_counter_4[103] <= 0;
        valid_bit_1[104]  <=   0;dirty_bit_1[104] <= 0;tag_address_1[104] <= 0;cache_block_1[104] <= 0;lru_counter_1[104] <= 0;valid_bit_2[104]  <=   0;dirty_bit_2[104] <= 0;tag_address_2[104] <= 0;cache_block_2[104] <= 0;lru_counter_2[104] <= 0;valid_bit_3[104]  <=   0;dirty_bit_3[104] <= 0;tag_address_3[104] <= 0;cache_block_3[104] <= 0;lru_counter_3[104] <= 0;valid_bit_4[104]  <=   0;dirty_bit_4[104] <= 0;tag_address_4[104] <= 0;cache_block_4[104] <= 0;lru_counter_4[104] <= 0;
        valid_bit_1[105]  <=   0;dirty_bit_1[105] <= 0;tag_address_1[105] <= 0;cache_block_1[105] <= 0;lru_counter_1[105] <= 0;valid_bit_2[105]  <=   0;dirty_bit_2[105] <= 0;tag_address_2[105] <= 0;cache_block_2[105] <= 0;lru_counter_2[105] <= 0;valid_bit_3[105]  <=   0;dirty_bit_3[105] <= 0;tag_address_3[105] <= 0;cache_block_3[105] <= 0;lru_counter_3[105] <= 0;valid_bit_4[105]  <=   0;dirty_bit_4[105] <= 0;tag_address_4[105] <= 0;cache_block_4[105] <= 0;lru_counter_4[105] <= 0;
        valid_bit_1[106]  <=   0;dirty_bit_1[106] <= 0;tag_address_1[106] <= 0;cache_block_1[106] <= 0;lru_counter_1[106] <= 0;valid_bit_2[106]  <=   0;dirty_bit_2[106] <= 0;tag_address_2[106] <= 0;cache_block_2[106] <= 0;lru_counter_2[106] <= 0;valid_bit_3[106]  <=   0;dirty_bit_3[106] <= 0;tag_address_3[106] <= 0;cache_block_3[106] <= 0;lru_counter_3[106] <= 0;valid_bit_4[106]  <=   0;dirty_bit_4[106] <= 0;tag_address_4[106] <= 0;cache_block_4[106] <= 0;lru_counter_4[106] <= 0;
        valid_bit_1[107]  <=   0;dirty_bit_1[107] <= 0;tag_address_1[107] <= 0;cache_block_1[107] <= 0;lru_counter_1[107] <= 0;valid_bit_2[107]  <=   0;dirty_bit_2[107] <= 0;tag_address_2[107] <= 0;cache_block_2[107] <= 0;lru_counter_2[107] <= 0;valid_bit_3[107]  <=   0;dirty_bit_3[107] <= 0;tag_address_3[107] <= 0;cache_block_3[107] <= 0;lru_counter_3[107] <= 0;valid_bit_4[107]  <=   0;dirty_bit_4[107] <= 0;tag_address_4[107] <= 0;cache_block_4[107] <= 0;lru_counter_4[107] <= 0;
        valid_bit_1[108]  <=   0;dirty_bit_1[108] <= 0;tag_address_1[108] <= 0;cache_block_1[108] <= 0;lru_counter_1[108] <= 0;valid_bit_2[108]  <=   0;dirty_bit_2[108] <= 0;tag_address_2[108] <= 0;cache_block_2[108] <= 0;lru_counter_2[108] <= 0;valid_bit_3[108]  <=   0;dirty_bit_3[108] <= 0;tag_address_3[108] <= 0;cache_block_3[108] <= 0;lru_counter_3[108] <= 0;valid_bit_4[108]  <=   0;dirty_bit_4[108] <= 0;tag_address_4[108] <= 0;cache_block_4[108] <= 0;lru_counter_4[108] <= 0;
        valid_bit_1[109]  <=   0;dirty_bit_1[109] <= 0;tag_address_1[109] <= 0;cache_block_1[109] <= 0;lru_counter_1[109] <= 0;valid_bit_2[109]  <=   0;dirty_bit_2[109] <= 0;tag_address_2[109] <= 0;cache_block_2[109] <= 0;lru_counter_2[109] <= 0;valid_bit_3[109]  <=   0;dirty_bit_3[109] <= 0;tag_address_3[109] <= 0;cache_block_3[109] <= 0;lru_counter_3[109] <= 0;valid_bit_4[109]  <=   0;dirty_bit_4[109] <= 0;tag_address_4[109] <= 0;cache_block_4[109] <= 0;lru_counter_4[109] <= 0;
        valid_bit_1[110]  <=   0;dirty_bit_1[110] <= 0;tag_address_1[110] <= 0;cache_block_1[110] <= 0;lru_counter_1[110] <= 0;valid_bit_2[110]  <=   0;dirty_bit_2[110] <= 0;tag_address_2[110] <= 0;cache_block_2[110] <= 0;lru_counter_2[110] <= 0;valid_bit_3[110]  <=   0;dirty_bit_3[110] <= 0;tag_address_3[110] <= 0;cache_block_3[110] <= 0;lru_counter_3[110] <= 0;valid_bit_4[110]  <=   0;dirty_bit_4[110] <= 0;tag_address_4[110] <= 0;cache_block_4[110] <= 0;lru_counter_4[110] <= 0;
        valid_bit_1[111]  <=   0;dirty_bit_1[111] <= 0;tag_address_1[111] <= 0;cache_block_1[111] <= 0;lru_counter_1[111] <= 0;valid_bit_2[111]  <=   0;dirty_bit_2[111] <= 0;tag_address_2[111] <= 0;cache_block_2[111] <= 0;lru_counter_2[111] <= 0;valid_bit_3[111]  <=   0;dirty_bit_3[111] <= 0;tag_address_3[111] <= 0;cache_block_3[111] <= 0;lru_counter_3[111] <= 0;valid_bit_4[111]  <=   0;dirty_bit_4[111] <= 0;tag_address_4[111] <= 0;cache_block_4[111] <= 0;lru_counter_4[111] <= 0;
        valid_bit_1[112]  <=   0;dirty_bit_1[112] <= 0;tag_address_1[112] <= 0;cache_block_1[112] <= 0;lru_counter_1[112] <= 0;valid_bit_2[112]  <=   0;dirty_bit_2[112] <= 0;tag_address_2[112] <= 0;cache_block_2[112] <= 0;lru_counter_2[112] <= 0;valid_bit_3[112]  <=   0;dirty_bit_3[112] <= 0;tag_address_3[112] <= 0;cache_block_3[112] <= 0;lru_counter_3[112] <= 0;valid_bit_4[112]  <=   0;dirty_bit_4[112] <= 0;tag_address_4[112] <= 0;cache_block_4[112] <= 0;lru_counter_4[112] <= 0;
        valid_bit_1[113]  <=   0;dirty_bit_1[113] <= 0;tag_address_1[113] <= 0;cache_block_1[113] <= 0;lru_counter_1[113] <= 0;valid_bit_2[113]  <=   0;dirty_bit_2[113] <= 0;tag_address_2[113] <= 0;cache_block_2[113] <= 0;lru_counter_2[113] <= 0;valid_bit_3[113]  <=   0;dirty_bit_3[113] <= 0;tag_address_3[113] <= 0;cache_block_3[113] <= 0;lru_counter_3[113] <= 0;valid_bit_4[113]  <=   0;dirty_bit_4[113] <= 0;tag_address_4[113] <= 0;cache_block_4[113] <= 0;lru_counter_4[113] <= 0;
        valid_bit_1[114]  <=   0;dirty_bit_1[114] <= 0;tag_address_1[114] <= 0;cache_block_1[114] <= 0;lru_counter_1[114] <= 0;valid_bit_2[114]  <=   0;dirty_bit_2[114] <= 0;tag_address_2[114] <= 0;cache_block_2[114] <= 0;lru_counter_2[114] <= 0;valid_bit_3[114]  <=   0;dirty_bit_3[114] <= 0;tag_address_3[114] <= 0;cache_block_3[114] <= 0;lru_counter_3[114] <= 0;valid_bit_4[114]  <=   0;dirty_bit_4[114] <= 0;tag_address_4[114] <= 0;cache_block_4[114] <= 0;lru_counter_4[114] <= 0;
        valid_bit_1[115]  <=   0;dirty_bit_1[115] <= 0;tag_address_1[115] <= 0;cache_block_1[115] <= 0;lru_counter_1[115] <= 0;valid_bit_2[115]  <=   0;dirty_bit_2[115] <= 0;tag_address_2[115] <= 0;cache_block_2[115] <= 0;lru_counter_2[115] <= 0;valid_bit_3[115]  <=   0;dirty_bit_3[115] <= 0;tag_address_3[115] <= 0;cache_block_3[115] <= 0;lru_counter_3[115] <= 0;valid_bit_4[115]  <=   0;dirty_bit_4[115] <= 0;tag_address_4[115] <= 0;cache_block_4[115] <= 0;lru_counter_4[115] <= 0;
        valid_bit_1[116]  <=   0;dirty_bit_1[116] <= 0;tag_address_1[116] <= 0;cache_block_1[116] <= 0;lru_counter_1[116] <= 0;valid_bit_2[116]  <=   0;dirty_bit_2[116] <= 0;tag_address_2[116] <= 0;cache_block_2[116] <= 0;lru_counter_2[116] <= 0;valid_bit_3[116]  <=   0;dirty_bit_3[116] <= 0;tag_address_3[116] <= 0;cache_block_3[116] <= 0;lru_counter_3[116] <= 0;valid_bit_4[116]  <=   0;dirty_bit_4[116] <= 0;tag_address_4[116] <= 0;cache_block_4[116] <= 0;lru_counter_4[116] <= 0;
        valid_bit_1[117]  <=   0;dirty_bit_1[117] <= 0;tag_address_1[117] <= 0;cache_block_1[117] <= 0;lru_counter_1[117] <= 0;valid_bit_2[117]  <=   0;dirty_bit_2[117] <= 0;tag_address_2[117] <= 0;cache_block_2[117] <= 0;lru_counter_2[117] <= 0;valid_bit_3[117]  <=   0;dirty_bit_3[117] <= 0;tag_address_3[117] <= 0;cache_block_3[117] <= 0;lru_counter_3[117] <= 0;valid_bit_4[117]  <=   0;dirty_bit_4[117] <= 0;tag_address_4[117] <= 0;cache_block_4[117] <= 0;lru_counter_4[117] <= 0;
        valid_bit_1[118]  <=   0;dirty_bit_1[118] <= 0;tag_address_1[118] <= 0;cache_block_1[118] <= 0;lru_counter_1[118] <= 0;valid_bit_2[118]  <=   0;dirty_bit_2[118] <= 0;tag_address_2[118] <= 0;cache_block_2[118] <= 0;lru_counter_2[118] <= 0;valid_bit_3[118]  <=   0;dirty_bit_3[118] <= 0;tag_address_3[118] <= 0;cache_block_3[118] <= 0;lru_counter_3[118] <= 0;valid_bit_4[118]  <=   0;dirty_bit_4[118] <= 0;tag_address_4[118] <= 0;cache_block_4[118] <= 0;lru_counter_4[118] <= 0;
        valid_bit_1[119]  <=   0;dirty_bit_1[119] <= 0;tag_address_1[119] <= 0;cache_block_1[119] <= 0;lru_counter_1[119] <= 0;valid_bit_2[119]  <=   0;dirty_bit_2[119] <= 0;tag_address_2[119] <= 0;cache_block_2[119] <= 0;lru_counter_2[119] <= 0;valid_bit_3[119]  <=   0;dirty_bit_3[119] <= 0;tag_address_3[119] <= 0;cache_block_3[119] <= 0;lru_counter_3[119] <= 0;valid_bit_4[119]  <=   0;dirty_bit_4[119] <= 0;tag_address_4[119] <= 0;cache_block_4[119] <= 0;lru_counter_4[119] <= 0;
        valid_bit_1[120]  <=   0;dirty_bit_1[120] <= 0;tag_address_1[120] <= 0;cache_block_1[120] <= 0;lru_counter_1[120] <= 0;valid_bit_2[120]  <=   0;dirty_bit_2[120] <= 0;tag_address_2[120] <= 0;cache_block_2[120] <= 0;lru_counter_2[120] <= 0;valid_bit_3[120]  <=   0;dirty_bit_3[120] <= 0;tag_address_3[120] <= 0;cache_block_3[120] <= 0;lru_counter_3[120] <= 0;valid_bit_4[120]  <=   0;dirty_bit_4[120] <= 0;tag_address_4[120] <= 0;cache_block_4[120] <= 0;lru_counter_4[120] <= 0;
        valid_bit_1[121]  <=   0;dirty_bit_1[121] <= 0;tag_address_1[121] <= 0;cache_block_1[121] <= 0;lru_counter_1[121] <= 0;valid_bit_2[121]  <=   0;dirty_bit_2[121] <= 0;tag_address_2[121] <= 0;cache_block_2[121] <= 0;lru_counter_2[121] <= 0;valid_bit_3[121]  <=   0;dirty_bit_3[121] <= 0;tag_address_3[121] <= 0;cache_block_3[121] <= 0;lru_counter_3[121] <= 0;valid_bit_4[121]  <=   0;dirty_bit_4[121] <= 0;tag_address_4[121] <= 0;cache_block_4[121] <= 0;lru_counter_4[121] <= 0;
        valid_bit_1[122]  <=   0;dirty_bit_1[122] <= 0;tag_address_1[122] <= 0;cache_block_1[122] <= 0;lru_counter_1[122] <= 0;valid_bit_2[122]  <=   0;dirty_bit_2[122] <= 0;tag_address_2[122] <= 0;cache_block_2[122] <= 0;lru_counter_2[122] <= 0;valid_bit_3[122]  <=   0;dirty_bit_3[122] <= 0;tag_address_3[122] <= 0;cache_block_3[122] <= 0;lru_counter_3[122] <= 0;valid_bit_4[122]  <=   0;dirty_bit_4[122] <= 0;tag_address_4[122] <= 0;cache_block_4[122] <= 0;lru_counter_4[122] <= 0;
        valid_bit_1[123]  <=   0;dirty_bit_1[123] <= 0;tag_address_1[123] <= 0;cache_block_1[123] <= 0;lru_counter_1[123] <= 0;valid_bit_2[123]  <=   0;dirty_bit_2[123] <= 0;tag_address_2[123] <= 0;cache_block_2[123] <= 0;lru_counter_2[123] <= 0;valid_bit_3[123]  <=   0;dirty_bit_3[123] <= 0;tag_address_3[123] <= 0;cache_block_3[123] <= 0;lru_counter_3[123] <= 0;valid_bit_4[123]  <=   0;dirty_bit_4[123] <= 0;tag_address_4[123] <= 0;cache_block_4[123] <= 0;lru_counter_4[123] <= 0;
        valid_bit_1[124]  <=   0;dirty_bit_1[124] <= 0;tag_address_1[124] <= 0;cache_block_1[124] <= 0;lru_counter_1[124] <= 0;valid_bit_2[124]  <=   0;dirty_bit_2[124] <= 0;tag_address_2[124] <= 0;cache_block_2[124] <= 0;lru_counter_2[124] <= 0;valid_bit_3[124]  <=   0;dirty_bit_3[124] <= 0;tag_address_3[124] <= 0;cache_block_3[124] <= 0;lru_counter_3[124] <= 0;valid_bit_4[124]  <=   0;dirty_bit_4[124] <= 0;tag_address_4[124] <= 0;cache_block_4[124] <= 0;lru_counter_4[124] <= 0;
        valid_bit_1[125]  <=   0;dirty_bit_1[125] <= 0;tag_address_1[125] <= 0;cache_block_1[125] <= 0;lru_counter_1[125] <= 0;valid_bit_2[125]  <=   0;dirty_bit_2[125] <= 0;tag_address_2[125] <= 0;cache_block_2[125] <= 0;lru_counter_2[125] <= 0;valid_bit_3[125]  <=   0;dirty_bit_3[125] <= 0;tag_address_3[125] <= 0;cache_block_3[125] <= 0;lru_counter_3[125] <= 0;valid_bit_4[125]  <=   0;dirty_bit_4[125] <= 0;tag_address_4[125] <= 0;cache_block_4[125] <= 0;lru_counter_4[125] <= 0;
        valid_bit_1[126]  <=   0;dirty_bit_1[126] <= 0;tag_address_1[126] <= 0;cache_block_1[126] <= 0;lru_counter_1[126] <= 0;valid_bit_2[126]  <=   0;dirty_bit_2[126] <= 0;tag_address_2[126] <= 0;cache_block_2[126] <= 0;lru_counter_2[126] <= 0;valid_bit_3[126]  <=   0;dirty_bit_3[126] <= 0;tag_address_3[126] <= 0;cache_block_3[126] <= 0;lru_counter_3[126] <= 0;valid_bit_4[126]  <=   0;dirty_bit_4[126] <= 0;tag_address_4[126] <= 0;cache_block_4[126] <= 0;lru_counter_4[126] <= 0;
        valid_bit_1[127]  <=   0;dirty_bit_1[127] <= 0;tag_address_1[127] <= 0;cache_block_1[127] <= 0;lru_counter_1[127] <= 0;valid_bit_2[127]  <=   0;dirty_bit_2[127] <= 0;tag_address_2[127] <= 0;cache_block_2[127] <= 0;lru_counter_2[127] <= 0;valid_bit_3[127]  <=   0;dirty_bit_3[127] <= 0;tag_address_3[127] <= 0;cache_block_3[127] <= 0;lru_counter_3[127] <= 0;valid_bit_4[127]  <=   0;dirty_bit_4[127] <= 0;tag_address_4[127] <= 0;cache_block_4[127] <= 0;lru_counter_4[127] <= 0;
        valid_bit_1[128]  <=   0;dirty_bit_1[128] <= 0;tag_address_1[128] <= 0;cache_block_1[128] <= 0;lru_counter_1[128] <= 0;valid_bit_2[128]  <=   0;dirty_bit_2[128] <= 0;tag_address_2[128] <= 0;cache_block_2[128] <= 0;lru_counter_2[128] <= 0;valid_bit_3[128]  <=   0;dirty_bit_3[128] <= 0;tag_address_3[128] <= 0;cache_block_3[128] <= 0;lru_counter_3[128] <= 0;valid_bit_4[128]  <=   0;dirty_bit_4[128] <= 0;tag_address_4[128] <= 0;cache_block_4[128] <= 0;lru_counter_4[128] <= 0;
        valid_bit_1[129]  <=   0;dirty_bit_1[129] <= 0;tag_address_1[129] <= 0;cache_block_1[129] <= 0;lru_counter_1[129] <= 0;valid_bit_2[129]  <=   0;dirty_bit_2[129] <= 0;tag_address_2[129] <= 0;cache_block_2[129] <= 0;lru_counter_2[129] <= 0;valid_bit_3[129]  <=   0;dirty_bit_3[129] <= 0;tag_address_3[129] <= 0;cache_block_3[129] <= 0;lru_counter_3[129] <= 0;valid_bit_4[129]  <=   0;dirty_bit_4[129] <= 0;tag_address_4[129] <= 0;cache_block_4[129] <= 0;lru_counter_4[129] <= 0;
        valid_bit_1[130]  <=   0;dirty_bit_1[130] <= 0;tag_address_1[130] <= 0;cache_block_1[130] <= 0;lru_counter_1[130] <= 0;valid_bit_2[130]  <=   0;dirty_bit_2[130] <= 0;tag_address_2[130] <= 0;cache_block_2[130] <= 0;lru_counter_2[130] <= 0;valid_bit_3[130]  <=   0;dirty_bit_3[130] <= 0;tag_address_3[130] <= 0;cache_block_3[130] <= 0;lru_counter_3[130] <= 0;valid_bit_4[130]  <=   0;dirty_bit_4[130] <= 0;tag_address_4[130] <= 0;cache_block_4[130] <= 0;lru_counter_4[130] <= 0;
        valid_bit_1[131]  <=   0;dirty_bit_1[131] <= 0;tag_address_1[131] <= 0;cache_block_1[131] <= 0;lru_counter_1[131] <= 0;valid_bit_2[131]  <=   0;dirty_bit_2[131] <= 0;tag_address_2[131] <= 0;cache_block_2[131] <= 0;lru_counter_2[131] <= 0;valid_bit_3[131]  <=   0;dirty_bit_3[131] <= 0;tag_address_3[131] <= 0;cache_block_3[131] <= 0;lru_counter_3[131] <= 0;valid_bit_4[131]  <=   0;dirty_bit_4[131] <= 0;tag_address_4[131] <= 0;cache_block_4[131] <= 0;lru_counter_4[131] <= 0;
        valid_bit_1[132]  <=   0;dirty_bit_1[132] <= 0;tag_address_1[132] <= 0;cache_block_1[132] <= 0;lru_counter_1[132] <= 0;valid_bit_2[132]  <=   0;dirty_bit_2[132] <= 0;tag_address_2[132] <= 0;cache_block_2[132] <= 0;lru_counter_2[132] <= 0;valid_bit_3[132]  <=   0;dirty_bit_3[132] <= 0;tag_address_3[132] <= 0;cache_block_3[132] <= 0;lru_counter_3[132] <= 0;valid_bit_4[132]  <=   0;dirty_bit_4[132] <= 0;tag_address_4[132] <= 0;cache_block_4[132] <= 0;lru_counter_4[132] <= 0;
        valid_bit_1[133]  <=   0;dirty_bit_1[133] <= 0;tag_address_1[133] <= 0;cache_block_1[133] <= 0;lru_counter_1[133] <= 0;valid_bit_2[133]  <=   0;dirty_bit_2[133] <= 0;tag_address_2[133] <= 0;cache_block_2[133] <= 0;lru_counter_2[133] <= 0;valid_bit_3[133]  <=   0;dirty_bit_3[133] <= 0;tag_address_3[133] <= 0;cache_block_3[133] <= 0;lru_counter_3[133] <= 0;valid_bit_4[133]  <=   0;dirty_bit_4[133] <= 0;tag_address_4[133] <= 0;cache_block_4[133] <= 0;lru_counter_4[133] <= 0;
        valid_bit_1[134]  <=   0;dirty_bit_1[134] <= 0;tag_address_1[134] <= 0;cache_block_1[134] <= 0;lru_counter_1[134] <= 0;valid_bit_2[134]  <=   0;dirty_bit_2[134] <= 0;tag_address_2[134] <= 0;cache_block_2[134] <= 0;lru_counter_2[134] <= 0;valid_bit_3[134]  <=   0;dirty_bit_3[134] <= 0;tag_address_3[134] <= 0;cache_block_3[134] <= 0;lru_counter_3[134] <= 0;valid_bit_4[134]  <=   0;dirty_bit_4[134] <= 0;tag_address_4[134] <= 0;cache_block_4[134] <= 0;lru_counter_4[134] <= 0;
        valid_bit_1[135]  <=   0;dirty_bit_1[135] <= 0;tag_address_1[135] <= 0;cache_block_1[135] <= 0;lru_counter_1[135] <= 0;valid_bit_2[135]  <=   0;dirty_bit_2[135] <= 0;tag_address_2[135] <= 0;cache_block_2[135] <= 0;lru_counter_2[135] <= 0;valid_bit_3[135]  <=   0;dirty_bit_3[135] <= 0;tag_address_3[135] <= 0;cache_block_3[135] <= 0;lru_counter_3[135] <= 0;valid_bit_4[135]  <=   0;dirty_bit_4[135] <= 0;tag_address_4[135] <= 0;cache_block_4[135] <= 0;lru_counter_4[135] <= 0;
        valid_bit_1[136]  <=   0;dirty_bit_1[136] <= 0;tag_address_1[136] <= 0;cache_block_1[136] <= 0;lru_counter_1[136] <= 0;valid_bit_2[136]  <=   0;dirty_bit_2[136] <= 0;tag_address_2[136] <= 0;cache_block_2[136] <= 0;lru_counter_2[136] <= 0;valid_bit_3[136]  <=   0;dirty_bit_3[136] <= 0;tag_address_3[136] <= 0;cache_block_3[136] <= 0;lru_counter_3[136] <= 0;valid_bit_4[136]  <=   0;dirty_bit_4[136] <= 0;tag_address_4[136] <= 0;cache_block_4[136] <= 0;lru_counter_4[136] <= 0;
        valid_bit_1[137]  <=   0;dirty_bit_1[137] <= 0;tag_address_1[137] <= 0;cache_block_1[137] <= 0;lru_counter_1[137] <= 0;valid_bit_2[137]  <=   0;dirty_bit_2[137] <= 0;tag_address_2[137] <= 0;cache_block_2[137] <= 0;lru_counter_2[137] <= 0;valid_bit_3[137]  <=   0;dirty_bit_3[137] <= 0;tag_address_3[137] <= 0;cache_block_3[137] <= 0;lru_counter_3[137] <= 0;valid_bit_4[137]  <=   0;dirty_bit_4[137] <= 0;tag_address_4[137] <= 0;cache_block_4[137] <= 0;lru_counter_4[137] <= 0;
        valid_bit_1[138]  <=   0;dirty_bit_1[138] <= 0;tag_address_1[138] <= 0;cache_block_1[138] <= 0;lru_counter_1[138] <= 0;valid_bit_2[138]  <=   0;dirty_bit_2[138] <= 0;tag_address_2[138] <= 0;cache_block_2[138] <= 0;lru_counter_2[138] <= 0;valid_bit_3[138]  <=   0;dirty_bit_3[138] <= 0;tag_address_3[138] <= 0;cache_block_3[138] <= 0;lru_counter_3[138] <= 0;valid_bit_4[138]  <=   0;dirty_bit_4[138] <= 0;tag_address_4[138] <= 0;cache_block_4[138] <= 0;lru_counter_4[138] <= 0;
        valid_bit_1[139]  <=   0;dirty_bit_1[139] <= 0;tag_address_1[139] <= 0;cache_block_1[139] <= 0;lru_counter_1[139] <= 0;valid_bit_2[139]  <=   0;dirty_bit_2[139] <= 0;tag_address_2[139] <= 0;cache_block_2[139] <= 0;lru_counter_2[139] <= 0;valid_bit_3[139]  <=   0;dirty_bit_3[139] <= 0;tag_address_3[139] <= 0;cache_block_3[139] <= 0;lru_counter_3[139] <= 0;valid_bit_4[139]  <=   0;dirty_bit_4[139] <= 0;tag_address_4[139] <= 0;cache_block_4[139] <= 0;lru_counter_4[139] <= 0;
        valid_bit_1[140]  <=   0;dirty_bit_1[140] <= 0;tag_address_1[140] <= 0;cache_block_1[140] <= 0;lru_counter_1[140] <= 0;valid_bit_2[140]  <=   0;dirty_bit_2[140] <= 0;tag_address_2[140] <= 0;cache_block_2[140] <= 0;lru_counter_2[140] <= 0;valid_bit_3[140]  <=   0;dirty_bit_3[140] <= 0;tag_address_3[140] <= 0;cache_block_3[140] <= 0;lru_counter_3[140] <= 0;valid_bit_4[140]  <=   0;dirty_bit_4[140] <= 0;tag_address_4[140] <= 0;cache_block_4[140] <= 0;lru_counter_4[140] <= 0;
        valid_bit_1[141]  <=   0;dirty_bit_1[141] <= 0;tag_address_1[141] <= 0;cache_block_1[141] <= 0;lru_counter_1[141] <= 0;valid_bit_2[141]  <=   0;dirty_bit_2[141] <= 0;tag_address_2[141] <= 0;cache_block_2[141] <= 0;lru_counter_2[141] <= 0;valid_bit_3[141]  <=   0;dirty_bit_3[141] <= 0;tag_address_3[141] <= 0;cache_block_3[141] <= 0;lru_counter_3[141] <= 0;valid_bit_4[141]  <=   0;dirty_bit_4[141] <= 0;tag_address_4[141] <= 0;cache_block_4[141] <= 0;lru_counter_4[141] <= 0;
        valid_bit_1[142]  <=   0;dirty_bit_1[142] <= 0;tag_address_1[142] <= 0;cache_block_1[142] <= 0;lru_counter_1[142] <= 0;valid_bit_2[142]  <=   0;dirty_bit_2[142] <= 0;tag_address_2[142] <= 0;cache_block_2[142] <= 0;lru_counter_2[142] <= 0;valid_bit_3[142]  <=   0;dirty_bit_3[142] <= 0;tag_address_3[142] <= 0;cache_block_3[142] <= 0;lru_counter_3[142] <= 0;valid_bit_4[142]  <=   0;dirty_bit_4[142] <= 0;tag_address_4[142] <= 0;cache_block_4[142] <= 0;lru_counter_4[142] <= 0;
        valid_bit_1[143]  <=   0;dirty_bit_1[143] <= 0;tag_address_1[143] <= 0;cache_block_1[143] <= 0;lru_counter_1[143] <= 0;valid_bit_2[143]  <=   0;dirty_bit_2[143] <= 0;tag_address_2[143] <= 0;cache_block_2[143] <= 0;lru_counter_2[143] <= 0;valid_bit_3[143]  <=   0;dirty_bit_3[143] <= 0;tag_address_3[143] <= 0;cache_block_3[143] <= 0;lru_counter_3[143] <= 0;valid_bit_4[143]  <=   0;dirty_bit_4[143] <= 0;tag_address_4[143] <= 0;cache_block_4[143] <= 0;lru_counter_4[143] <= 0;
        valid_bit_1[144]  <=   0;dirty_bit_1[144] <= 0;tag_address_1[144] <= 0;cache_block_1[144] <= 0;lru_counter_1[144] <= 0;valid_bit_2[144]  <=   0;dirty_bit_2[144] <= 0;tag_address_2[144] <= 0;cache_block_2[144] <= 0;lru_counter_2[144] <= 0;valid_bit_3[144]  <=   0;dirty_bit_3[144] <= 0;tag_address_3[144] <= 0;cache_block_3[144] <= 0;lru_counter_3[144] <= 0;valid_bit_4[144]  <=   0;dirty_bit_4[144] <= 0;tag_address_4[144] <= 0;cache_block_4[144] <= 0;lru_counter_4[144] <= 0;
        valid_bit_1[145]  <=   0;dirty_bit_1[145] <= 0;tag_address_1[145] <= 0;cache_block_1[145] <= 0;lru_counter_1[145] <= 0;valid_bit_2[145]  <=   0;dirty_bit_2[145] <= 0;tag_address_2[145] <= 0;cache_block_2[145] <= 0;lru_counter_2[145] <= 0;valid_bit_3[145]  <=   0;dirty_bit_3[145] <= 0;tag_address_3[145] <= 0;cache_block_3[145] <= 0;lru_counter_3[145] <= 0;valid_bit_4[145]  <=   0;dirty_bit_4[145] <= 0;tag_address_4[145] <= 0;cache_block_4[145] <= 0;lru_counter_4[145] <= 0;
        valid_bit_1[146]  <=   0;dirty_bit_1[146] <= 0;tag_address_1[146] <= 0;cache_block_1[146] <= 0;lru_counter_1[146] <= 0;valid_bit_2[146]  <=   0;dirty_bit_2[146] <= 0;tag_address_2[146] <= 0;cache_block_2[146] <= 0;lru_counter_2[146] <= 0;valid_bit_3[146]  <=   0;dirty_bit_3[146] <= 0;tag_address_3[146] <= 0;cache_block_3[146] <= 0;lru_counter_3[146] <= 0;valid_bit_4[146]  <=   0;dirty_bit_4[146] <= 0;tag_address_4[146] <= 0;cache_block_4[146] <= 0;lru_counter_4[146] <= 0;
        valid_bit_1[147]  <=   0;dirty_bit_1[147] <= 0;tag_address_1[147] <= 0;cache_block_1[147] <= 0;lru_counter_1[147] <= 0;valid_bit_2[147]  <=   0;dirty_bit_2[147] <= 0;tag_address_2[147] <= 0;cache_block_2[147] <= 0;lru_counter_2[147] <= 0;valid_bit_3[147]  <=   0;dirty_bit_3[147] <= 0;tag_address_3[147] <= 0;cache_block_3[147] <= 0;lru_counter_3[147] <= 0;valid_bit_4[147]  <=   0;dirty_bit_4[147] <= 0;tag_address_4[147] <= 0;cache_block_4[147] <= 0;lru_counter_4[147] <= 0;
        valid_bit_1[148]  <=   0;dirty_bit_1[148] <= 0;tag_address_1[148] <= 0;cache_block_1[148] <= 0;lru_counter_1[148] <= 0;valid_bit_2[148]  <=   0;dirty_bit_2[148] <= 0;tag_address_2[148] <= 0;cache_block_2[148] <= 0;lru_counter_2[148] <= 0;valid_bit_3[148]  <=   0;dirty_bit_3[148] <= 0;tag_address_3[148] <= 0;cache_block_3[148] <= 0;lru_counter_3[148] <= 0;valid_bit_4[148]  <=   0;dirty_bit_4[148] <= 0;tag_address_4[148] <= 0;cache_block_4[148] <= 0;lru_counter_4[148] <= 0;
        valid_bit_1[149]  <=   0;dirty_bit_1[149] <= 0;tag_address_1[149] <= 0;cache_block_1[149] <= 0;lru_counter_1[149] <= 0;valid_bit_2[149]  <=   0;dirty_bit_2[149] <= 0;tag_address_2[149] <= 0;cache_block_2[149] <= 0;lru_counter_2[149] <= 0;valid_bit_3[149]  <=   0;dirty_bit_3[149] <= 0;tag_address_3[149] <= 0;cache_block_3[149] <= 0;lru_counter_3[149] <= 0;valid_bit_4[149]  <=   0;dirty_bit_4[149] <= 0;tag_address_4[149] <= 0;cache_block_4[149] <= 0;lru_counter_4[149] <= 0;
        valid_bit_1[150]  <=   0;dirty_bit_1[150] <= 0;tag_address_1[150] <= 0;cache_block_1[150] <= 0;lru_counter_1[150] <= 0;valid_bit_2[150]  <=   0;dirty_bit_2[150] <= 0;tag_address_2[150] <= 0;cache_block_2[150] <= 0;lru_counter_2[150] <= 0;valid_bit_3[150]  <=   0;dirty_bit_3[150] <= 0;tag_address_3[150] <= 0;cache_block_3[150] <= 0;lru_counter_3[150] <= 0;valid_bit_4[150]  <=   0;dirty_bit_4[150] <= 0;tag_address_4[150] <= 0;cache_block_4[150] <= 0;lru_counter_4[150] <= 0;
        valid_bit_1[151]  <=   0;dirty_bit_1[151] <= 0;tag_address_1[151] <= 0;cache_block_1[151] <= 0;lru_counter_1[151] <= 0;valid_bit_2[151]  <=   0;dirty_bit_2[151] <= 0;tag_address_2[151] <= 0;cache_block_2[151] <= 0;lru_counter_2[151] <= 0;valid_bit_3[151]  <=   0;dirty_bit_3[151] <= 0;tag_address_3[151] <= 0;cache_block_3[151] <= 0;lru_counter_3[151] <= 0;valid_bit_4[151]  <=   0;dirty_bit_4[151] <= 0;tag_address_4[151] <= 0;cache_block_4[151] <= 0;lru_counter_4[151] <= 0;
        valid_bit_1[152]  <=   0;dirty_bit_1[152] <= 0;tag_address_1[152] <= 0;cache_block_1[152] <= 0;lru_counter_1[152] <= 0;valid_bit_2[152]  <=   0;dirty_bit_2[152] <= 0;tag_address_2[152] <= 0;cache_block_2[152] <= 0;lru_counter_2[152] <= 0;valid_bit_3[152]  <=   0;dirty_bit_3[152] <= 0;tag_address_3[152] <= 0;cache_block_3[152] <= 0;lru_counter_3[152] <= 0;valid_bit_4[152]  <=   0;dirty_bit_4[152] <= 0;tag_address_4[152] <= 0;cache_block_4[152] <= 0;lru_counter_4[152] <= 0;
        valid_bit_1[153]  <=   0;dirty_bit_1[153] <= 0;tag_address_1[153] <= 0;cache_block_1[153] <= 0;lru_counter_1[153] <= 0;valid_bit_2[153]  <=   0;dirty_bit_2[153] <= 0;tag_address_2[153] <= 0;cache_block_2[153] <= 0;lru_counter_2[153] <= 0;valid_bit_3[153]  <=   0;dirty_bit_3[153] <= 0;tag_address_3[153] <= 0;cache_block_3[153] <= 0;lru_counter_3[153] <= 0;valid_bit_4[153]  <=   0;dirty_bit_4[153] <= 0;tag_address_4[153] <= 0;cache_block_4[153] <= 0;lru_counter_4[153] <= 0;
        valid_bit_1[154]  <=   0;dirty_bit_1[154] <= 0;tag_address_1[154] <= 0;cache_block_1[154] <= 0;lru_counter_1[154] <= 0;valid_bit_2[154]  <=   0;dirty_bit_2[154] <= 0;tag_address_2[154] <= 0;cache_block_2[154] <= 0;lru_counter_2[154] <= 0;valid_bit_3[154]  <=   0;dirty_bit_3[154] <= 0;tag_address_3[154] <= 0;cache_block_3[154] <= 0;lru_counter_3[154] <= 0;valid_bit_4[154]  <=   0;dirty_bit_4[154] <= 0;tag_address_4[154] <= 0;cache_block_4[154] <= 0;lru_counter_4[154] <= 0;
        valid_bit_1[155]  <=   0;dirty_bit_1[155] <= 0;tag_address_1[155] <= 0;cache_block_1[155] <= 0;lru_counter_1[155] <= 0;valid_bit_2[155]  <=   0;dirty_bit_2[155] <= 0;tag_address_2[155] <= 0;cache_block_2[155] <= 0;lru_counter_2[155] <= 0;valid_bit_3[155]  <=   0;dirty_bit_3[155] <= 0;tag_address_3[155] <= 0;cache_block_3[155] <= 0;lru_counter_3[155] <= 0;valid_bit_4[155]  <=   0;dirty_bit_4[155] <= 0;tag_address_4[155] <= 0;cache_block_4[155] <= 0;lru_counter_4[155] <= 0;
        valid_bit_1[156]  <=   0;dirty_bit_1[156] <= 0;tag_address_1[156] <= 0;cache_block_1[156] <= 0;lru_counter_1[156] <= 0;valid_bit_2[156]  <=   0;dirty_bit_2[156] <= 0;tag_address_2[156] <= 0;cache_block_2[156] <= 0;lru_counter_2[156] <= 0;valid_bit_3[156]  <=   0;dirty_bit_3[156] <= 0;tag_address_3[156] <= 0;cache_block_3[156] <= 0;lru_counter_3[156] <= 0;valid_bit_4[156]  <=   0;dirty_bit_4[156] <= 0;tag_address_4[156] <= 0;cache_block_4[156] <= 0;lru_counter_4[156] <= 0;
        valid_bit_1[157]  <=   0;dirty_bit_1[157] <= 0;tag_address_1[157] <= 0;cache_block_1[157] <= 0;lru_counter_1[157] <= 0;valid_bit_2[157]  <=   0;dirty_bit_2[157] <= 0;tag_address_2[157] <= 0;cache_block_2[157] <= 0;lru_counter_2[157] <= 0;valid_bit_3[157]  <=   0;dirty_bit_3[157] <= 0;tag_address_3[157] <= 0;cache_block_3[157] <= 0;lru_counter_3[157] <= 0;valid_bit_4[157]  <=   0;dirty_bit_4[157] <= 0;tag_address_4[157] <= 0;cache_block_4[157] <= 0;lru_counter_4[157] <= 0;
        valid_bit_1[158]  <=   0;dirty_bit_1[158] <= 0;tag_address_1[158] <= 0;cache_block_1[158] <= 0;lru_counter_1[158] <= 0;valid_bit_2[158]  <=   0;dirty_bit_2[158] <= 0;tag_address_2[158] <= 0;cache_block_2[158] <= 0;lru_counter_2[158] <= 0;valid_bit_3[158]  <=   0;dirty_bit_3[158] <= 0;tag_address_3[158] <= 0;cache_block_3[158] <= 0;lru_counter_3[158] <= 0;valid_bit_4[158]  <=   0;dirty_bit_4[158] <= 0;tag_address_4[158] <= 0;cache_block_4[158] <= 0;lru_counter_4[158] <= 0;
        valid_bit_1[159]  <=   0;dirty_bit_1[159] <= 0;tag_address_1[159] <= 0;cache_block_1[159] <= 0;lru_counter_1[159] <= 0;valid_bit_2[159]  <=   0;dirty_bit_2[159] <= 0;tag_address_2[159] <= 0;cache_block_2[159] <= 0;lru_counter_2[159] <= 0;valid_bit_3[159]  <=   0;dirty_bit_3[159] <= 0;tag_address_3[159] <= 0;cache_block_3[159] <= 0;lru_counter_3[159] <= 0;valid_bit_4[159]  <=   0;dirty_bit_4[159] <= 0;tag_address_4[159] <= 0;cache_block_4[159] <= 0;lru_counter_4[159] <= 0;
        valid_bit_1[160]  <=   0;dirty_bit_1[160] <= 0;tag_address_1[160] <= 0;cache_block_1[160] <= 0;lru_counter_1[160] <= 0;valid_bit_2[160]  <=   0;dirty_bit_2[160] <= 0;tag_address_2[160] <= 0;cache_block_2[160] <= 0;lru_counter_2[160] <= 0;valid_bit_3[160]  <=   0;dirty_bit_3[160] <= 0;tag_address_3[160] <= 0;cache_block_3[160] <= 0;lru_counter_3[160] <= 0;valid_bit_4[160]  <=   0;dirty_bit_4[160] <= 0;tag_address_4[160] <= 0;cache_block_4[160] <= 0;lru_counter_4[160] <= 0;
        valid_bit_1[161]  <=   0;dirty_bit_1[161] <= 0;tag_address_1[161] <= 0;cache_block_1[161] <= 0;lru_counter_1[161] <= 0;valid_bit_2[161]  <=   0;dirty_bit_2[161] <= 0;tag_address_2[161] <= 0;cache_block_2[161] <= 0;lru_counter_2[161] <= 0;valid_bit_3[161]  <=   0;dirty_bit_3[161] <= 0;tag_address_3[161] <= 0;cache_block_3[161] <= 0;lru_counter_3[161] <= 0;valid_bit_4[161]  <=   0;dirty_bit_4[161] <= 0;tag_address_4[161] <= 0;cache_block_4[161] <= 0;lru_counter_4[161] <= 0;
        valid_bit_1[162]  <=   0;dirty_bit_1[162] <= 0;tag_address_1[162] <= 0;cache_block_1[162] <= 0;lru_counter_1[162] <= 0;valid_bit_2[162]  <=   0;dirty_bit_2[162] <= 0;tag_address_2[162] <= 0;cache_block_2[162] <= 0;lru_counter_2[162] <= 0;valid_bit_3[162]  <=   0;dirty_bit_3[162] <= 0;tag_address_3[162] <= 0;cache_block_3[162] <= 0;lru_counter_3[162] <= 0;valid_bit_4[162]  <=   0;dirty_bit_4[162] <= 0;tag_address_4[162] <= 0;cache_block_4[162] <= 0;lru_counter_4[162] <= 0;
        valid_bit_1[163]  <=   0;dirty_bit_1[163] <= 0;tag_address_1[163] <= 0;cache_block_1[163] <= 0;lru_counter_1[163] <= 0;valid_bit_2[163]  <=   0;dirty_bit_2[163] <= 0;tag_address_2[163] <= 0;cache_block_2[163] <= 0;lru_counter_2[163] <= 0;valid_bit_3[163]  <=   0;dirty_bit_3[163] <= 0;tag_address_3[163] <= 0;cache_block_3[163] <= 0;lru_counter_3[163] <= 0;valid_bit_4[163]  <=   0;dirty_bit_4[163] <= 0;tag_address_4[163] <= 0;cache_block_4[163] <= 0;lru_counter_4[163] <= 0;
        valid_bit_1[164]  <=   0;dirty_bit_1[164] <= 0;tag_address_1[164] <= 0;cache_block_1[164] <= 0;lru_counter_1[164] <= 0;valid_bit_2[164]  <=   0;dirty_bit_2[164] <= 0;tag_address_2[164] <= 0;cache_block_2[164] <= 0;lru_counter_2[164] <= 0;valid_bit_3[164]  <=   0;dirty_bit_3[164] <= 0;tag_address_3[164] <= 0;cache_block_3[164] <= 0;lru_counter_3[164] <= 0;valid_bit_4[164]  <=   0;dirty_bit_4[164] <= 0;tag_address_4[164] <= 0;cache_block_4[164] <= 0;lru_counter_4[164] <= 0;
        valid_bit_1[165]  <=   0;dirty_bit_1[165] <= 0;tag_address_1[165] <= 0;cache_block_1[165] <= 0;lru_counter_1[165] <= 0;valid_bit_2[165]  <=   0;dirty_bit_2[165] <= 0;tag_address_2[165] <= 0;cache_block_2[165] <= 0;lru_counter_2[165] <= 0;valid_bit_3[165]  <=   0;dirty_bit_3[165] <= 0;tag_address_3[165] <= 0;cache_block_3[165] <= 0;lru_counter_3[165] <= 0;valid_bit_4[165]  <=   0;dirty_bit_4[165] <= 0;tag_address_4[165] <= 0;cache_block_4[165] <= 0;lru_counter_4[165] <= 0;
        valid_bit_1[166]  <=   0;dirty_bit_1[166] <= 0;tag_address_1[166] <= 0;cache_block_1[166] <= 0;lru_counter_1[166] <= 0;valid_bit_2[166]  <=   0;dirty_bit_2[166] <= 0;tag_address_2[166] <= 0;cache_block_2[166] <= 0;lru_counter_2[166] <= 0;valid_bit_3[166]  <=   0;dirty_bit_3[166] <= 0;tag_address_3[166] <= 0;cache_block_3[166] <= 0;lru_counter_3[166] <= 0;valid_bit_4[166]  <=   0;dirty_bit_4[166] <= 0;tag_address_4[166] <= 0;cache_block_4[166] <= 0;lru_counter_4[166] <= 0;
        valid_bit_1[167]  <=   0;dirty_bit_1[167] <= 0;tag_address_1[167] <= 0;cache_block_1[167] <= 0;lru_counter_1[167] <= 0;valid_bit_2[167]  <=   0;dirty_bit_2[167] <= 0;tag_address_2[167] <= 0;cache_block_2[167] <= 0;lru_counter_2[167] <= 0;valid_bit_3[167]  <=   0;dirty_bit_3[167] <= 0;tag_address_3[167] <= 0;cache_block_3[167] <= 0;lru_counter_3[167] <= 0;valid_bit_4[167]  <=   0;dirty_bit_4[167] <= 0;tag_address_4[167] <= 0;cache_block_4[167] <= 0;lru_counter_4[167] <= 0;
        valid_bit_1[168]  <=   0;dirty_bit_1[168] <= 0;tag_address_1[168] <= 0;cache_block_1[168] <= 0;lru_counter_1[168] <= 0;valid_bit_2[168]  <=   0;dirty_bit_2[168] <= 0;tag_address_2[168] <= 0;cache_block_2[168] <= 0;lru_counter_2[168] <= 0;valid_bit_3[168]  <=   0;dirty_bit_3[168] <= 0;tag_address_3[168] <= 0;cache_block_3[168] <= 0;lru_counter_3[168] <= 0;valid_bit_4[168]  <=   0;dirty_bit_4[168] <= 0;tag_address_4[168] <= 0;cache_block_4[168] <= 0;lru_counter_4[168] <= 0;
        valid_bit_1[169]  <=   0;dirty_bit_1[169] <= 0;tag_address_1[169] <= 0;cache_block_1[169] <= 0;lru_counter_1[169] <= 0;valid_bit_2[169]  <=   0;dirty_bit_2[169] <= 0;tag_address_2[169] <= 0;cache_block_2[169] <= 0;lru_counter_2[169] <= 0;valid_bit_3[169]  <=   0;dirty_bit_3[169] <= 0;tag_address_3[169] <= 0;cache_block_3[169] <= 0;lru_counter_3[169] <= 0;valid_bit_4[169]  <=   0;dirty_bit_4[169] <= 0;tag_address_4[169] <= 0;cache_block_4[169] <= 0;lru_counter_4[169] <= 0;
        valid_bit_1[170]  <=   0;dirty_bit_1[170] <= 0;tag_address_1[170] <= 0;cache_block_1[170] <= 0;lru_counter_1[170] <= 0;valid_bit_2[170]  <=   0;dirty_bit_2[170] <= 0;tag_address_2[170] <= 0;cache_block_2[170] <= 0;lru_counter_2[170] <= 0;valid_bit_3[170]  <=   0;dirty_bit_3[170] <= 0;tag_address_3[170] <= 0;cache_block_3[170] <= 0;lru_counter_3[170] <= 0;valid_bit_4[170]  <=   0;dirty_bit_4[170] <= 0;tag_address_4[170] <= 0;cache_block_4[170] <= 0;lru_counter_4[170] <= 0;
        valid_bit_1[171]  <=   0;dirty_bit_1[171] <= 0;tag_address_1[171] <= 0;cache_block_1[171] <= 0;lru_counter_1[171] <= 0;valid_bit_2[171]  <=   0;dirty_bit_2[171] <= 0;tag_address_2[171] <= 0;cache_block_2[171] <= 0;lru_counter_2[171] <= 0;valid_bit_3[171]  <=   0;dirty_bit_3[171] <= 0;tag_address_3[171] <= 0;cache_block_3[171] <= 0;lru_counter_3[171] <= 0;valid_bit_4[171]  <=   0;dirty_bit_4[171] <= 0;tag_address_4[171] <= 0;cache_block_4[171] <= 0;lru_counter_4[171] <= 0;
        valid_bit_1[172]  <=   0;dirty_bit_1[172] <= 0;tag_address_1[172] <= 0;cache_block_1[172] <= 0;lru_counter_1[172] <= 0;valid_bit_2[172]  <=   0;dirty_bit_2[172] <= 0;tag_address_2[172] <= 0;cache_block_2[172] <= 0;lru_counter_2[172] <= 0;valid_bit_3[172]  <=   0;dirty_bit_3[172] <= 0;tag_address_3[172] <= 0;cache_block_3[172] <= 0;lru_counter_3[172] <= 0;valid_bit_4[172]  <=   0;dirty_bit_4[172] <= 0;tag_address_4[172] <= 0;cache_block_4[172] <= 0;lru_counter_4[172] <= 0;
        valid_bit_1[173]  <=   0;dirty_bit_1[173] <= 0;tag_address_1[173] <= 0;cache_block_1[173] <= 0;lru_counter_1[173] <= 0;valid_bit_2[173]  <=   0;dirty_bit_2[173] <= 0;tag_address_2[173] <= 0;cache_block_2[173] <= 0;lru_counter_2[173] <= 0;valid_bit_3[173]  <=   0;dirty_bit_3[173] <= 0;tag_address_3[173] <= 0;cache_block_3[173] <= 0;lru_counter_3[173] <= 0;valid_bit_4[173]  <=   0;dirty_bit_4[173] <= 0;tag_address_4[173] <= 0;cache_block_4[173] <= 0;lru_counter_4[173] <= 0;
        valid_bit_1[174]  <=   0;dirty_bit_1[174] <= 0;tag_address_1[174] <= 0;cache_block_1[174] <= 0;lru_counter_1[174] <= 0;valid_bit_2[174]  <=   0;dirty_bit_2[174] <= 0;tag_address_2[174] <= 0;cache_block_2[174] <= 0;lru_counter_2[174] <= 0;valid_bit_3[174]  <=   0;dirty_bit_3[174] <= 0;tag_address_3[174] <= 0;cache_block_3[174] <= 0;lru_counter_3[174] <= 0;valid_bit_4[174]  <=   0;dirty_bit_4[174] <= 0;tag_address_4[174] <= 0;cache_block_4[174] <= 0;lru_counter_4[174] <= 0;
        valid_bit_1[175]  <=   0;dirty_bit_1[175] <= 0;tag_address_1[175] <= 0;cache_block_1[175] <= 0;lru_counter_1[175] <= 0;valid_bit_2[175]  <=   0;dirty_bit_2[175] <= 0;tag_address_2[175] <= 0;cache_block_2[175] <= 0;lru_counter_2[175] <= 0;valid_bit_3[175]  <=   0;dirty_bit_3[175] <= 0;tag_address_3[175] <= 0;cache_block_3[175] <= 0;lru_counter_3[175] <= 0;valid_bit_4[175]  <=   0;dirty_bit_4[175] <= 0;tag_address_4[175] <= 0;cache_block_4[175] <= 0;lru_counter_4[175] <= 0;
        valid_bit_1[176]  <=   0;dirty_bit_1[176] <= 0;tag_address_1[176] <= 0;cache_block_1[176] <= 0;lru_counter_1[176] <= 0;valid_bit_2[176]  <=   0;dirty_bit_2[176] <= 0;tag_address_2[176] <= 0;cache_block_2[176] <= 0;lru_counter_2[176] <= 0;valid_bit_3[176]  <=   0;dirty_bit_3[176] <= 0;tag_address_3[176] <= 0;cache_block_3[176] <= 0;lru_counter_3[176] <= 0;valid_bit_4[176]  <=   0;dirty_bit_4[176] <= 0;tag_address_4[176] <= 0;cache_block_4[176] <= 0;lru_counter_4[176] <= 0;
        valid_bit_1[177]  <=   0;dirty_bit_1[177] <= 0;tag_address_1[177] <= 0;cache_block_1[177] <= 0;lru_counter_1[177] <= 0;valid_bit_2[177]  <=   0;dirty_bit_2[177] <= 0;tag_address_2[177] <= 0;cache_block_2[177] <= 0;lru_counter_2[177] <= 0;valid_bit_3[177]  <=   0;dirty_bit_3[177] <= 0;tag_address_3[177] <= 0;cache_block_3[177] <= 0;lru_counter_3[177] <= 0;valid_bit_4[177]  <=   0;dirty_bit_4[177] <= 0;tag_address_4[177] <= 0;cache_block_4[177] <= 0;lru_counter_4[177] <= 0;
        valid_bit_1[178]  <=   0;dirty_bit_1[178] <= 0;tag_address_1[178] <= 0;cache_block_1[178] <= 0;lru_counter_1[178] <= 0;valid_bit_2[178]  <=   0;dirty_bit_2[178] <= 0;tag_address_2[178] <= 0;cache_block_2[178] <= 0;lru_counter_2[178] <= 0;valid_bit_3[178]  <=   0;dirty_bit_3[178] <= 0;tag_address_3[178] <= 0;cache_block_3[178] <= 0;lru_counter_3[178] <= 0;valid_bit_4[178]  <=   0;dirty_bit_4[178] <= 0;tag_address_4[178] <= 0;cache_block_4[178] <= 0;lru_counter_4[178] <= 0;
        valid_bit_1[179]  <=   0;dirty_bit_1[179] <= 0;tag_address_1[179] <= 0;cache_block_1[179] <= 0;lru_counter_1[179] <= 0;valid_bit_2[179]  <=   0;dirty_bit_2[179] <= 0;tag_address_2[179] <= 0;cache_block_2[179] <= 0;lru_counter_2[179] <= 0;valid_bit_3[179]  <=   0;dirty_bit_3[179] <= 0;tag_address_3[179] <= 0;cache_block_3[179] <= 0;lru_counter_3[179] <= 0;valid_bit_4[179]  <=   0;dirty_bit_4[179] <= 0;tag_address_4[179] <= 0;cache_block_4[179] <= 0;lru_counter_4[179] <= 0;
        valid_bit_1[180]  <=   0;dirty_bit_1[180] <= 0;tag_address_1[180] <= 0;cache_block_1[180] <= 0;lru_counter_1[180] <= 0;valid_bit_2[180]  <=   0;dirty_bit_2[180] <= 0;tag_address_2[180] <= 0;cache_block_2[180] <= 0;lru_counter_2[180] <= 0;valid_bit_3[180]  <=   0;dirty_bit_3[180] <= 0;tag_address_3[180] <= 0;cache_block_3[180] <= 0;lru_counter_3[180] <= 0;valid_bit_4[180]  <=   0;dirty_bit_4[180] <= 0;tag_address_4[180] <= 0;cache_block_4[180] <= 0;lru_counter_4[180] <= 0;
        valid_bit_1[181]  <=   0;dirty_bit_1[181] <= 0;tag_address_1[181] <= 0;cache_block_1[181] <= 0;lru_counter_1[181] <= 0;valid_bit_2[181]  <=   0;dirty_bit_2[181] <= 0;tag_address_2[181] <= 0;cache_block_2[181] <= 0;lru_counter_2[181] <= 0;valid_bit_3[181]  <=   0;dirty_bit_3[181] <= 0;tag_address_3[181] <= 0;cache_block_3[181] <= 0;lru_counter_3[181] <= 0;valid_bit_4[181]  <=   0;dirty_bit_4[181] <= 0;tag_address_4[181] <= 0;cache_block_4[181] <= 0;lru_counter_4[181] <= 0;
        valid_bit_1[182]  <=   0;dirty_bit_1[182] <= 0;tag_address_1[182] <= 0;cache_block_1[182] <= 0;lru_counter_1[182] <= 0;valid_bit_2[182]  <=   0;dirty_bit_2[182] <= 0;tag_address_2[182] <= 0;cache_block_2[182] <= 0;lru_counter_2[182] <= 0;valid_bit_3[182]  <=   0;dirty_bit_3[182] <= 0;tag_address_3[182] <= 0;cache_block_3[182] <= 0;lru_counter_3[182] <= 0;valid_bit_4[182]  <=   0;dirty_bit_4[182] <= 0;tag_address_4[182] <= 0;cache_block_4[182] <= 0;lru_counter_4[182] <= 0;
        valid_bit_1[183]  <=   0;dirty_bit_1[183] <= 0;tag_address_1[183] <= 0;cache_block_1[183] <= 0;lru_counter_1[183] <= 0;valid_bit_2[183]  <=   0;dirty_bit_2[183] <= 0;tag_address_2[183] <= 0;cache_block_2[183] <= 0;lru_counter_2[183] <= 0;valid_bit_3[183]  <=   0;dirty_bit_3[183] <= 0;tag_address_3[183] <= 0;cache_block_3[183] <= 0;lru_counter_3[183] <= 0;valid_bit_4[183]  <=   0;dirty_bit_4[183] <= 0;tag_address_4[183] <= 0;cache_block_4[183] <= 0;lru_counter_4[183] <= 0;
        valid_bit_1[184]  <=   0;dirty_bit_1[184] <= 0;tag_address_1[184] <= 0;cache_block_1[184] <= 0;lru_counter_1[184] <= 0;valid_bit_2[184]  <=   0;dirty_bit_2[184] <= 0;tag_address_2[184] <= 0;cache_block_2[184] <= 0;lru_counter_2[184] <= 0;valid_bit_3[184]  <=   0;dirty_bit_3[184] <= 0;tag_address_3[184] <= 0;cache_block_3[184] <= 0;lru_counter_3[184] <= 0;valid_bit_4[184]  <=   0;dirty_bit_4[184] <= 0;tag_address_4[184] <= 0;cache_block_4[184] <= 0;lru_counter_4[184] <= 0;
        valid_bit_1[185]  <=   0;dirty_bit_1[185] <= 0;tag_address_1[185] <= 0;cache_block_1[185] <= 0;lru_counter_1[185] <= 0;valid_bit_2[185]  <=   0;dirty_bit_2[185] <= 0;tag_address_2[185] <= 0;cache_block_2[185] <= 0;lru_counter_2[185] <= 0;valid_bit_3[185]  <=   0;dirty_bit_3[185] <= 0;tag_address_3[185] <= 0;cache_block_3[185] <= 0;lru_counter_3[185] <= 0;valid_bit_4[185]  <=   0;dirty_bit_4[185] <= 0;tag_address_4[185] <= 0;cache_block_4[185] <= 0;lru_counter_4[185] <= 0;
        valid_bit_1[186]  <=   0;dirty_bit_1[186] <= 0;tag_address_1[186] <= 0;cache_block_1[186] <= 0;lru_counter_1[186] <= 0;valid_bit_2[186]  <=   0;dirty_bit_2[186] <= 0;tag_address_2[186] <= 0;cache_block_2[186] <= 0;lru_counter_2[186] <= 0;valid_bit_3[186]  <=   0;dirty_bit_3[186] <= 0;tag_address_3[186] <= 0;cache_block_3[186] <= 0;lru_counter_3[186] <= 0;valid_bit_4[186]  <=   0;dirty_bit_4[186] <= 0;tag_address_4[186] <= 0;cache_block_4[186] <= 0;lru_counter_4[186] <= 0;
        valid_bit_1[187]  <=   0;dirty_bit_1[187] <= 0;tag_address_1[187] <= 0;cache_block_1[187] <= 0;lru_counter_1[187] <= 0;valid_bit_2[187]  <=   0;dirty_bit_2[187] <= 0;tag_address_2[187] <= 0;cache_block_2[187] <= 0;lru_counter_2[187] <= 0;valid_bit_3[187]  <=   0;dirty_bit_3[187] <= 0;tag_address_3[187] <= 0;cache_block_3[187] <= 0;lru_counter_3[187] <= 0;valid_bit_4[187]  <=   0;dirty_bit_4[187] <= 0;tag_address_4[187] <= 0;cache_block_4[187] <= 0;lru_counter_4[187] <= 0;
        valid_bit_1[188]  <=   0;dirty_bit_1[188] <= 0;tag_address_1[188] <= 0;cache_block_1[188] <= 0;lru_counter_1[188] <= 0;valid_bit_2[188]  <=   0;dirty_bit_2[188] <= 0;tag_address_2[188] <= 0;cache_block_2[188] <= 0;lru_counter_2[188] <= 0;valid_bit_3[188]  <=   0;dirty_bit_3[188] <= 0;tag_address_3[188] <= 0;cache_block_3[188] <= 0;lru_counter_3[188] <= 0;valid_bit_4[188]  <=   0;dirty_bit_4[188] <= 0;tag_address_4[188] <= 0;cache_block_4[188] <= 0;lru_counter_4[188] <= 0;
        valid_bit_1[189]  <=   0;dirty_bit_1[189] <= 0;tag_address_1[189] <= 0;cache_block_1[189] <= 0;lru_counter_1[189] <= 0;valid_bit_2[189]  <=   0;dirty_bit_2[189] <= 0;tag_address_2[189] <= 0;cache_block_2[189] <= 0;lru_counter_2[189] <= 0;valid_bit_3[189]  <=   0;dirty_bit_3[189] <= 0;tag_address_3[189] <= 0;cache_block_3[189] <= 0;lru_counter_3[189] <= 0;valid_bit_4[189]  <=   0;dirty_bit_4[189] <= 0;tag_address_4[189] <= 0;cache_block_4[189] <= 0;lru_counter_4[189] <= 0;
        valid_bit_1[190]  <=   0;dirty_bit_1[190] <= 0;tag_address_1[190] <= 0;cache_block_1[190] <= 0;lru_counter_1[190] <= 0;valid_bit_2[190]  <=   0;dirty_bit_2[190] <= 0;tag_address_2[190] <= 0;cache_block_2[190] <= 0;lru_counter_2[190] <= 0;valid_bit_3[190]  <=   0;dirty_bit_3[190] <= 0;tag_address_3[190] <= 0;cache_block_3[190] <= 0;lru_counter_3[190] <= 0;valid_bit_4[190]  <=   0;dirty_bit_4[190] <= 0;tag_address_4[190] <= 0;cache_block_4[190] <= 0;lru_counter_4[190] <= 0;
        valid_bit_1[191]  <=   0;dirty_bit_1[191] <= 0;tag_address_1[191] <= 0;cache_block_1[191] <= 0;lru_counter_1[191] <= 0;valid_bit_2[191]  <=   0;dirty_bit_2[191] <= 0;tag_address_2[191] <= 0;cache_block_2[191] <= 0;lru_counter_2[191] <= 0;valid_bit_3[191]  <=   0;dirty_bit_3[191] <= 0;tag_address_3[191] <= 0;cache_block_3[191] <= 0;lru_counter_3[191] <= 0;valid_bit_4[191]  <=   0;dirty_bit_4[191] <= 0;tag_address_4[191] <= 0;cache_block_4[191] <= 0;lru_counter_4[191] <= 0;
        valid_bit_1[192]  <=   0;dirty_bit_1[192] <= 0;tag_address_1[192] <= 0;cache_block_1[192] <= 0;lru_counter_1[192] <= 0;valid_bit_2[192]  <=   0;dirty_bit_2[192] <= 0;tag_address_2[192] <= 0;cache_block_2[192] <= 0;lru_counter_2[192] <= 0;valid_bit_3[192]  <=   0;dirty_bit_3[192] <= 0;tag_address_3[192] <= 0;cache_block_3[192] <= 0;lru_counter_3[192] <= 0;valid_bit_4[192]  <=   0;dirty_bit_4[192] <= 0;tag_address_4[192] <= 0;cache_block_4[192] <= 0;lru_counter_4[192] <= 0;
        valid_bit_1[193]  <=   0;dirty_bit_1[193] <= 0;tag_address_1[193] <= 0;cache_block_1[193] <= 0;lru_counter_1[193] <= 0;valid_bit_2[193]  <=   0;dirty_bit_2[193] <= 0;tag_address_2[193] <= 0;cache_block_2[193] <= 0;lru_counter_2[193] <= 0;valid_bit_3[193]  <=   0;dirty_bit_3[193] <= 0;tag_address_3[193] <= 0;cache_block_3[193] <= 0;lru_counter_3[193] <= 0;valid_bit_4[193]  <=   0;dirty_bit_4[193] <= 0;tag_address_4[193] <= 0;cache_block_4[193] <= 0;lru_counter_4[193] <= 0;
        valid_bit_1[194]  <=   0;dirty_bit_1[194] <= 0;tag_address_1[194] <= 0;cache_block_1[194] <= 0;lru_counter_1[194] <= 0;valid_bit_2[194]  <=   0;dirty_bit_2[194] <= 0;tag_address_2[194] <= 0;cache_block_2[194] <= 0;lru_counter_2[194] <= 0;valid_bit_3[194]  <=   0;dirty_bit_3[194] <= 0;tag_address_3[194] <= 0;cache_block_3[194] <= 0;lru_counter_3[194] <= 0;valid_bit_4[194]  <=   0;dirty_bit_4[194] <= 0;tag_address_4[194] <= 0;cache_block_4[194] <= 0;lru_counter_4[194] <= 0;
        valid_bit_1[195]  <=   0;dirty_bit_1[195] <= 0;tag_address_1[195] <= 0;cache_block_1[195] <= 0;lru_counter_1[195] <= 0;valid_bit_2[195]  <=   0;dirty_bit_2[195] <= 0;tag_address_2[195] <= 0;cache_block_2[195] <= 0;lru_counter_2[195] <= 0;valid_bit_3[195]  <=   0;dirty_bit_3[195] <= 0;tag_address_3[195] <= 0;cache_block_3[195] <= 0;lru_counter_3[195] <= 0;valid_bit_4[195]  <=   0;dirty_bit_4[195] <= 0;tag_address_4[195] <= 0;cache_block_4[195] <= 0;lru_counter_4[195] <= 0;
        valid_bit_1[196]  <=   0;dirty_bit_1[196] <= 0;tag_address_1[196] <= 0;cache_block_1[196] <= 0;lru_counter_1[196] <= 0;valid_bit_2[196]  <=   0;dirty_bit_2[196] <= 0;tag_address_2[196] <= 0;cache_block_2[196] <= 0;lru_counter_2[196] <= 0;valid_bit_3[196]  <=   0;dirty_bit_3[196] <= 0;tag_address_3[196] <= 0;cache_block_3[196] <= 0;lru_counter_3[196] <= 0;valid_bit_4[196]  <=   0;dirty_bit_4[196] <= 0;tag_address_4[196] <= 0;cache_block_4[196] <= 0;lru_counter_4[196] <= 0;
        valid_bit_1[197]  <=   0;dirty_bit_1[197] <= 0;tag_address_1[197] <= 0;cache_block_1[197] <= 0;lru_counter_1[197] <= 0;valid_bit_2[197]  <=   0;dirty_bit_2[197] <= 0;tag_address_2[197] <= 0;cache_block_2[197] <= 0;lru_counter_2[197] <= 0;valid_bit_3[197]  <=   0;dirty_bit_3[197] <= 0;tag_address_3[197] <= 0;cache_block_3[197] <= 0;lru_counter_3[197] <= 0;valid_bit_4[197]  <=   0;dirty_bit_4[197] <= 0;tag_address_4[197] <= 0;cache_block_4[197] <= 0;lru_counter_4[197] <= 0;
        valid_bit_1[198]  <=   0;dirty_bit_1[198] <= 0;tag_address_1[198] <= 0;cache_block_1[198] <= 0;lru_counter_1[198] <= 0;valid_bit_2[198]  <=   0;dirty_bit_2[198] <= 0;tag_address_2[198] <= 0;cache_block_2[198] <= 0;lru_counter_2[198] <= 0;valid_bit_3[198]  <=   0;dirty_bit_3[198] <= 0;tag_address_3[198] <= 0;cache_block_3[198] <= 0;lru_counter_3[198] <= 0;valid_bit_4[198]  <=   0;dirty_bit_4[198] <= 0;tag_address_4[198] <= 0;cache_block_4[198] <= 0;lru_counter_4[198] <= 0;
        valid_bit_1[199]  <=   0;dirty_bit_1[199] <= 0;tag_address_1[199] <= 0;cache_block_1[199] <= 0;lru_counter_1[199] <= 0;valid_bit_2[199]  <=   0;dirty_bit_2[199] <= 0;tag_address_2[199] <= 0;cache_block_2[199] <= 0;lru_counter_2[199] <= 0;valid_bit_3[199]  <=   0;dirty_bit_3[199] <= 0;tag_address_3[199] <= 0;cache_block_3[199] <= 0;lru_counter_3[199] <= 0;valid_bit_4[199]  <=   0;dirty_bit_4[199] <= 0;tag_address_4[199] <= 0;cache_block_4[199] <= 0;lru_counter_4[199] <= 0;
        valid_bit_1[200]  <=   0;dirty_bit_1[200] <= 0;tag_address_1[200] <= 0;cache_block_1[200] <= 0;lru_counter_1[200] <= 0;valid_bit_2[200]  <=   0;dirty_bit_2[200] <= 0;tag_address_2[200] <= 0;cache_block_2[200] <= 0;lru_counter_2[200] <= 0;valid_bit_3[200]  <=   0;dirty_bit_3[200] <= 0;tag_address_3[200] <= 0;cache_block_3[200] <= 0;lru_counter_3[200] <= 0;valid_bit_4[200]  <=   0;dirty_bit_4[200] <= 0;tag_address_4[200] <= 0;cache_block_4[200] <= 0;lru_counter_4[200] <= 0;
        valid_bit_1[201]  <=   0;dirty_bit_1[201] <= 0;tag_address_1[201] <= 0;cache_block_1[201] <= 0;lru_counter_1[201] <= 0;valid_bit_2[201]  <=   0;dirty_bit_2[201] <= 0;tag_address_2[201] <= 0;cache_block_2[201] <= 0;lru_counter_2[201] <= 0;valid_bit_3[201]  <=   0;dirty_bit_3[201] <= 0;tag_address_3[201] <= 0;cache_block_3[201] <= 0;lru_counter_3[201] <= 0;valid_bit_4[201]  <=   0;dirty_bit_4[201] <= 0;tag_address_4[201] <= 0;cache_block_4[201] <= 0;lru_counter_4[201] <= 0;
        valid_bit_1[202]  <=   0;dirty_bit_1[202] <= 0;tag_address_1[202] <= 0;cache_block_1[202] <= 0;lru_counter_1[202] <= 0;valid_bit_2[202]  <=   0;dirty_bit_2[202] <= 0;tag_address_2[202] <= 0;cache_block_2[202] <= 0;lru_counter_2[202] <= 0;valid_bit_3[202]  <=   0;dirty_bit_3[202] <= 0;tag_address_3[202] <= 0;cache_block_3[202] <= 0;lru_counter_3[202] <= 0;valid_bit_4[202]  <=   0;dirty_bit_4[202] <= 0;tag_address_4[202] <= 0;cache_block_4[202] <= 0;lru_counter_4[202] <= 0;
        valid_bit_1[203]  <=   0;dirty_bit_1[203] <= 0;tag_address_1[203] <= 0;cache_block_1[203] <= 0;lru_counter_1[203] <= 0;valid_bit_2[203]  <=   0;dirty_bit_2[203] <= 0;tag_address_2[203] <= 0;cache_block_2[203] <= 0;lru_counter_2[203] <= 0;valid_bit_3[203]  <=   0;dirty_bit_3[203] <= 0;tag_address_3[203] <= 0;cache_block_3[203] <= 0;lru_counter_3[203] <= 0;valid_bit_4[203]  <=   0;dirty_bit_4[203] <= 0;tag_address_4[203] <= 0;cache_block_4[203] <= 0;lru_counter_4[203] <= 0;
        valid_bit_1[204]  <=   0;dirty_bit_1[204] <= 0;tag_address_1[204] <= 0;cache_block_1[204] <= 0;lru_counter_1[204] <= 0;valid_bit_2[204]  <=   0;dirty_bit_2[204] <= 0;tag_address_2[204] <= 0;cache_block_2[204] <= 0;lru_counter_2[204] <= 0;valid_bit_3[204]  <=   0;dirty_bit_3[204] <= 0;tag_address_3[204] <= 0;cache_block_3[204] <= 0;lru_counter_3[204] <= 0;valid_bit_4[204]  <=   0;dirty_bit_4[204] <= 0;tag_address_4[204] <= 0;cache_block_4[204] <= 0;lru_counter_4[204] <= 0;
        valid_bit_1[205]  <=   0;dirty_bit_1[205] <= 0;tag_address_1[205] <= 0;cache_block_1[205] <= 0;lru_counter_1[205] <= 0;valid_bit_2[205]  <=   0;dirty_bit_2[205] <= 0;tag_address_2[205] <= 0;cache_block_2[205] <= 0;lru_counter_2[205] <= 0;valid_bit_3[205]  <=   0;dirty_bit_3[205] <= 0;tag_address_3[205] <= 0;cache_block_3[205] <= 0;lru_counter_3[205] <= 0;valid_bit_4[205]  <=   0;dirty_bit_4[205] <= 0;tag_address_4[205] <= 0;cache_block_4[205] <= 0;lru_counter_4[205] <= 0;
        valid_bit_1[206]  <=   0;dirty_bit_1[206] <= 0;tag_address_1[206] <= 0;cache_block_1[206] <= 0;lru_counter_1[206] <= 0;valid_bit_2[206]  <=   0;dirty_bit_2[206] <= 0;tag_address_2[206] <= 0;cache_block_2[206] <= 0;lru_counter_2[206] <= 0;valid_bit_3[206]  <=   0;dirty_bit_3[206] <= 0;tag_address_3[206] <= 0;cache_block_3[206] <= 0;lru_counter_3[206] <= 0;valid_bit_4[206]  <=   0;dirty_bit_4[206] <= 0;tag_address_4[206] <= 0;cache_block_4[206] <= 0;lru_counter_4[206] <= 0;
        valid_bit_1[207]  <=   0;dirty_bit_1[207] <= 0;tag_address_1[207] <= 0;cache_block_1[207] <= 0;lru_counter_1[207] <= 0;valid_bit_2[207]  <=   0;dirty_bit_2[207] <= 0;tag_address_2[207] <= 0;cache_block_2[207] <= 0;lru_counter_2[207] <= 0;valid_bit_3[207]  <=   0;dirty_bit_3[207] <= 0;tag_address_3[207] <= 0;cache_block_3[207] <= 0;lru_counter_3[207] <= 0;valid_bit_4[207]  <=   0;dirty_bit_4[207] <= 0;tag_address_4[207] <= 0;cache_block_4[207] <= 0;lru_counter_4[207] <= 0;
        valid_bit_1[208]  <=   0;dirty_bit_1[208] <= 0;tag_address_1[208] <= 0;cache_block_1[208] <= 0;lru_counter_1[208] <= 0;valid_bit_2[208]  <=   0;dirty_bit_2[208] <= 0;tag_address_2[208] <= 0;cache_block_2[208] <= 0;lru_counter_2[208] <= 0;valid_bit_3[208]  <=   0;dirty_bit_3[208] <= 0;tag_address_3[208] <= 0;cache_block_3[208] <= 0;lru_counter_3[208] <= 0;valid_bit_4[208]  <=   0;dirty_bit_4[208] <= 0;tag_address_4[208] <= 0;cache_block_4[208] <= 0;lru_counter_4[208] <= 0;
        valid_bit_1[209]  <=   0;dirty_bit_1[209] <= 0;tag_address_1[209] <= 0;cache_block_1[209] <= 0;lru_counter_1[209] <= 0;valid_bit_2[209]  <=   0;dirty_bit_2[209] <= 0;tag_address_2[209] <= 0;cache_block_2[209] <= 0;lru_counter_2[209] <= 0;valid_bit_3[209]  <=   0;dirty_bit_3[209] <= 0;tag_address_3[209] <= 0;cache_block_3[209] <= 0;lru_counter_3[209] <= 0;valid_bit_4[209]  <=   0;dirty_bit_4[209] <= 0;tag_address_4[209] <= 0;cache_block_4[209] <= 0;lru_counter_4[209] <= 0;
        valid_bit_1[210]  <=   0;dirty_bit_1[210] <= 0;tag_address_1[210] <= 0;cache_block_1[210] <= 0;lru_counter_1[210] <= 0;valid_bit_2[210]  <=   0;dirty_bit_2[210] <= 0;tag_address_2[210] <= 0;cache_block_2[210] <= 0;lru_counter_2[210] <= 0;valid_bit_3[210]  <=   0;dirty_bit_3[210] <= 0;tag_address_3[210] <= 0;cache_block_3[210] <= 0;lru_counter_3[210] <= 0;valid_bit_4[210]  <=   0;dirty_bit_4[210] <= 0;tag_address_4[210] <= 0;cache_block_4[210] <= 0;lru_counter_4[210] <= 0;
        valid_bit_1[211]  <=   0;dirty_bit_1[211] <= 0;tag_address_1[211] <= 0;cache_block_1[211] <= 0;lru_counter_1[211] <= 0;valid_bit_2[211]  <=   0;dirty_bit_2[211] <= 0;tag_address_2[211] <= 0;cache_block_2[211] <= 0;lru_counter_2[211] <= 0;valid_bit_3[211]  <=   0;dirty_bit_3[211] <= 0;tag_address_3[211] <= 0;cache_block_3[211] <= 0;lru_counter_3[211] <= 0;valid_bit_4[211]  <=   0;dirty_bit_4[211] <= 0;tag_address_4[211] <= 0;cache_block_4[211] <= 0;lru_counter_4[211] <= 0;
        valid_bit_1[212]  <=   0;dirty_bit_1[212] <= 0;tag_address_1[212] <= 0;cache_block_1[212] <= 0;lru_counter_1[212] <= 0;valid_bit_2[212]  <=   0;dirty_bit_2[212] <= 0;tag_address_2[212] <= 0;cache_block_2[212] <= 0;lru_counter_2[212] <= 0;valid_bit_3[212]  <=   0;dirty_bit_3[212] <= 0;tag_address_3[212] <= 0;cache_block_3[212] <= 0;lru_counter_3[212] <= 0;valid_bit_4[212]  <=   0;dirty_bit_4[212] <= 0;tag_address_4[212] <= 0;cache_block_4[212] <= 0;lru_counter_4[212] <= 0;
        valid_bit_1[213]  <=   0;dirty_bit_1[213] <= 0;tag_address_1[213] <= 0;cache_block_1[213] <= 0;lru_counter_1[213] <= 0;valid_bit_2[213]  <=   0;dirty_bit_2[213] <= 0;tag_address_2[213] <= 0;cache_block_2[213] <= 0;lru_counter_2[213] <= 0;valid_bit_3[213]  <=   0;dirty_bit_3[213] <= 0;tag_address_3[213] <= 0;cache_block_3[213] <= 0;lru_counter_3[213] <= 0;valid_bit_4[213]  <=   0;dirty_bit_4[213] <= 0;tag_address_4[213] <= 0;cache_block_4[213] <= 0;lru_counter_4[213] <= 0;
        valid_bit_1[214]  <=   0;dirty_bit_1[214] <= 0;tag_address_1[214] <= 0;cache_block_1[214] <= 0;lru_counter_1[214] <= 0;valid_bit_2[214]  <=   0;dirty_bit_2[214] <= 0;tag_address_2[214] <= 0;cache_block_2[214] <= 0;lru_counter_2[214] <= 0;valid_bit_3[214]  <=   0;dirty_bit_3[214] <= 0;tag_address_3[214] <= 0;cache_block_3[214] <= 0;lru_counter_3[214] <= 0;valid_bit_4[214]  <=   0;dirty_bit_4[214] <= 0;tag_address_4[214] <= 0;cache_block_4[214] <= 0;lru_counter_4[214] <= 0;
        valid_bit_1[215]  <=   0;dirty_bit_1[215] <= 0;tag_address_1[215] <= 0;cache_block_1[215] <= 0;lru_counter_1[215] <= 0;valid_bit_2[215]  <=   0;dirty_bit_2[215] <= 0;tag_address_2[215] <= 0;cache_block_2[215] <= 0;lru_counter_2[215] <= 0;valid_bit_3[215]  <=   0;dirty_bit_3[215] <= 0;tag_address_3[215] <= 0;cache_block_3[215] <= 0;lru_counter_3[215] <= 0;valid_bit_4[215]  <=   0;dirty_bit_4[215] <= 0;tag_address_4[215] <= 0;cache_block_4[215] <= 0;lru_counter_4[215] <= 0;
        valid_bit_1[216]  <=   0;dirty_bit_1[216] <= 0;tag_address_1[216] <= 0;cache_block_1[216] <= 0;lru_counter_1[216] <= 0;valid_bit_2[216]  <=   0;dirty_bit_2[216] <= 0;tag_address_2[216] <= 0;cache_block_2[216] <= 0;lru_counter_2[216] <= 0;valid_bit_3[216]  <=   0;dirty_bit_3[216] <= 0;tag_address_3[216] <= 0;cache_block_3[216] <= 0;lru_counter_3[216] <= 0;valid_bit_4[216]  <=   0;dirty_bit_4[216] <= 0;tag_address_4[216] <= 0;cache_block_4[216] <= 0;lru_counter_4[216] <= 0;
        valid_bit_1[217]  <=   0;dirty_bit_1[217] <= 0;tag_address_1[217] <= 0;cache_block_1[217] <= 0;lru_counter_1[217] <= 0;valid_bit_2[217]  <=   0;dirty_bit_2[217] <= 0;tag_address_2[217] <= 0;cache_block_2[217] <= 0;lru_counter_2[217] <= 0;valid_bit_3[217]  <=   0;dirty_bit_3[217] <= 0;tag_address_3[217] <= 0;cache_block_3[217] <= 0;lru_counter_3[217] <= 0;valid_bit_4[217]  <=   0;dirty_bit_4[217] <= 0;tag_address_4[217] <= 0;cache_block_4[217] <= 0;lru_counter_4[217] <= 0;
        valid_bit_1[218]  <=   0;dirty_bit_1[218] <= 0;tag_address_1[218] <= 0;cache_block_1[218] <= 0;lru_counter_1[218] <= 0;valid_bit_2[218]  <=   0;dirty_bit_2[218] <= 0;tag_address_2[218] <= 0;cache_block_2[218] <= 0;lru_counter_2[218] <= 0;valid_bit_3[218]  <=   0;dirty_bit_3[218] <= 0;tag_address_3[218] <= 0;cache_block_3[218] <= 0;lru_counter_3[218] <= 0;valid_bit_4[218]  <=   0;dirty_bit_4[218] <= 0;tag_address_4[218] <= 0;cache_block_4[218] <= 0;lru_counter_4[218] <= 0;
        valid_bit_1[219]  <=   0;dirty_bit_1[219] <= 0;tag_address_1[219] <= 0;cache_block_1[219] <= 0;lru_counter_1[219] <= 0;valid_bit_2[219]  <=   0;dirty_bit_2[219] <= 0;tag_address_2[219] <= 0;cache_block_2[219] <= 0;lru_counter_2[219] <= 0;valid_bit_3[219]  <=   0;dirty_bit_3[219] <= 0;tag_address_3[219] <= 0;cache_block_3[219] <= 0;lru_counter_3[219] <= 0;valid_bit_4[219]  <=   0;dirty_bit_4[219] <= 0;tag_address_4[219] <= 0;cache_block_4[219] <= 0;lru_counter_4[219] <= 0;
        valid_bit_1[220]  <=   0;dirty_bit_1[220] <= 0;tag_address_1[220] <= 0;cache_block_1[220] <= 0;lru_counter_1[220] <= 0;valid_bit_2[220]  <=   0;dirty_bit_2[220] <= 0;tag_address_2[220] <= 0;cache_block_2[220] <= 0;lru_counter_2[220] <= 0;valid_bit_3[220]  <=   0;dirty_bit_3[220] <= 0;tag_address_3[220] <= 0;cache_block_3[220] <= 0;lru_counter_3[220] <= 0;valid_bit_4[220]  <=   0;dirty_bit_4[220] <= 0;tag_address_4[220] <= 0;cache_block_4[220] <= 0;lru_counter_4[220] <= 0;
        valid_bit_1[221]  <=   0;dirty_bit_1[221] <= 0;tag_address_1[221] <= 0;cache_block_1[221] <= 0;lru_counter_1[221] <= 0;valid_bit_2[221]  <=   0;dirty_bit_2[221] <= 0;tag_address_2[221] <= 0;cache_block_2[221] <= 0;lru_counter_2[221] <= 0;valid_bit_3[221]  <=   0;dirty_bit_3[221] <= 0;tag_address_3[221] <= 0;cache_block_3[221] <= 0;lru_counter_3[221] <= 0;valid_bit_4[221]  <=   0;dirty_bit_4[221] <= 0;tag_address_4[221] <= 0;cache_block_4[221] <= 0;lru_counter_4[221] <= 0;
        valid_bit_1[222]  <=   0;dirty_bit_1[222] <= 0;tag_address_1[222] <= 0;cache_block_1[222] <= 0;lru_counter_1[222] <= 0;valid_bit_2[222]  <=   0;dirty_bit_2[222] <= 0;tag_address_2[222] <= 0;cache_block_2[222] <= 0;lru_counter_2[222] <= 0;valid_bit_3[222]  <=   0;dirty_bit_3[222] <= 0;tag_address_3[222] <= 0;cache_block_3[222] <= 0;lru_counter_3[222] <= 0;valid_bit_4[222]  <=   0;dirty_bit_4[222] <= 0;tag_address_4[222] <= 0;cache_block_4[222] <= 0;lru_counter_4[222] <= 0;
        valid_bit_1[223]  <=   0;dirty_bit_1[223] <= 0;tag_address_1[223] <= 0;cache_block_1[223] <= 0;lru_counter_1[223] <= 0;valid_bit_2[223]  <=   0;dirty_bit_2[223] <= 0;tag_address_2[223] <= 0;cache_block_2[223] <= 0;lru_counter_2[223] <= 0;valid_bit_3[223]  <=   0;dirty_bit_3[223] <= 0;tag_address_3[223] <= 0;cache_block_3[223] <= 0;lru_counter_3[223] <= 0;valid_bit_4[223]  <=   0;dirty_bit_4[223] <= 0;tag_address_4[223] <= 0;cache_block_4[223] <= 0;lru_counter_4[223] <= 0;
        valid_bit_1[224]  <=   0;dirty_bit_1[224] <= 0;tag_address_1[224] <= 0;cache_block_1[224] <= 0;lru_counter_1[224] <= 0;valid_bit_2[224]  <=   0;dirty_bit_2[224] <= 0;tag_address_2[224] <= 0;cache_block_2[224] <= 0;lru_counter_2[224] <= 0;valid_bit_3[224]  <=   0;dirty_bit_3[224] <= 0;tag_address_3[224] <= 0;cache_block_3[224] <= 0;lru_counter_3[224] <= 0;valid_bit_4[224]  <=   0;dirty_bit_4[224] <= 0;tag_address_4[224] <= 0;cache_block_4[224] <= 0;lru_counter_4[224] <= 0;
        valid_bit_1[225]  <=   0;dirty_bit_1[225] <= 0;tag_address_1[225] <= 0;cache_block_1[225] <= 0;lru_counter_1[225] <= 0;valid_bit_2[225]  <=   0;dirty_bit_2[225] <= 0;tag_address_2[225] <= 0;cache_block_2[225] <= 0;lru_counter_2[225] <= 0;valid_bit_3[225]  <=   0;dirty_bit_3[225] <= 0;tag_address_3[225] <= 0;cache_block_3[225] <= 0;lru_counter_3[225] <= 0;valid_bit_4[225]  <=   0;dirty_bit_4[225] <= 0;tag_address_4[225] <= 0;cache_block_4[225] <= 0;lru_counter_4[225] <= 0;
        valid_bit_1[226]  <=   0;dirty_bit_1[226] <= 0;tag_address_1[226] <= 0;cache_block_1[226] <= 0;lru_counter_1[226] <= 0;valid_bit_2[226]  <=   0;dirty_bit_2[226] <= 0;tag_address_2[226] <= 0;cache_block_2[226] <= 0;lru_counter_2[226] <= 0;valid_bit_3[226]  <=   0;dirty_bit_3[226] <= 0;tag_address_3[226] <= 0;cache_block_3[226] <= 0;lru_counter_3[226] <= 0;valid_bit_4[226]  <=   0;dirty_bit_4[226] <= 0;tag_address_4[226] <= 0;cache_block_4[226] <= 0;lru_counter_4[226] <= 0;
        valid_bit_1[227]  <=   0;dirty_bit_1[227] <= 0;tag_address_1[227] <= 0;cache_block_1[227] <= 0;lru_counter_1[227] <= 0;valid_bit_2[227]  <=   0;dirty_bit_2[227] <= 0;tag_address_2[227] <= 0;cache_block_2[227] <= 0;lru_counter_2[227] <= 0;valid_bit_3[227]  <=   0;dirty_bit_3[227] <= 0;tag_address_3[227] <= 0;cache_block_3[227] <= 0;lru_counter_3[227] <= 0;valid_bit_4[227]  <=   0;dirty_bit_4[227] <= 0;tag_address_4[227] <= 0;cache_block_4[227] <= 0;lru_counter_4[227] <= 0;
        valid_bit_1[228]  <=   0;dirty_bit_1[228] <= 0;tag_address_1[228] <= 0;cache_block_1[228] <= 0;lru_counter_1[228] <= 0;valid_bit_2[228]  <=   0;dirty_bit_2[228] <= 0;tag_address_2[228] <= 0;cache_block_2[228] <= 0;lru_counter_2[228] <= 0;valid_bit_3[228]  <=   0;dirty_bit_3[228] <= 0;tag_address_3[228] <= 0;cache_block_3[228] <= 0;lru_counter_3[228] <= 0;valid_bit_4[228]  <=   0;dirty_bit_4[228] <= 0;tag_address_4[228] <= 0;cache_block_4[228] <= 0;lru_counter_4[228] <= 0;
        valid_bit_1[229]  <=   0;dirty_bit_1[229] <= 0;tag_address_1[229] <= 0;cache_block_1[229] <= 0;lru_counter_1[229] <= 0;valid_bit_2[229]  <=   0;dirty_bit_2[229] <= 0;tag_address_2[229] <= 0;cache_block_2[229] <= 0;lru_counter_2[229] <= 0;valid_bit_3[229]  <=   0;dirty_bit_3[229] <= 0;tag_address_3[229] <= 0;cache_block_3[229] <= 0;lru_counter_3[229] <= 0;valid_bit_4[229]  <=   0;dirty_bit_4[229] <= 0;tag_address_4[229] <= 0;cache_block_4[229] <= 0;lru_counter_4[229] <= 0;
        valid_bit_1[230]  <=   0;dirty_bit_1[230] <= 0;tag_address_1[230] <= 0;cache_block_1[230] <= 0;lru_counter_1[230] <= 0;valid_bit_2[230]  <=   0;dirty_bit_2[230] <= 0;tag_address_2[230] <= 0;cache_block_2[230] <= 0;lru_counter_2[230] <= 0;valid_bit_3[230]  <=   0;dirty_bit_3[230] <= 0;tag_address_3[230] <= 0;cache_block_3[230] <= 0;lru_counter_3[230] <= 0;valid_bit_4[230]  <=   0;dirty_bit_4[230] <= 0;tag_address_4[230] <= 0;cache_block_4[230] <= 0;lru_counter_4[230] <= 0;
        valid_bit_1[231]  <=   0;dirty_bit_1[231] <= 0;tag_address_1[231] <= 0;cache_block_1[231] <= 0;lru_counter_1[231] <= 0;valid_bit_2[231]  <=   0;dirty_bit_2[231] <= 0;tag_address_2[231] <= 0;cache_block_2[231] <= 0;lru_counter_2[231] <= 0;valid_bit_3[231]  <=   0;dirty_bit_3[231] <= 0;tag_address_3[231] <= 0;cache_block_3[231] <= 0;lru_counter_3[231] <= 0;valid_bit_4[231]  <=   0;dirty_bit_4[231] <= 0;tag_address_4[231] <= 0;cache_block_4[231] <= 0;lru_counter_4[231] <= 0;
        valid_bit_1[232]  <=   0;dirty_bit_1[232] <= 0;tag_address_1[232] <= 0;cache_block_1[232] <= 0;lru_counter_1[232] <= 0;valid_bit_2[232]  <=   0;dirty_bit_2[232] <= 0;tag_address_2[232] <= 0;cache_block_2[232] <= 0;lru_counter_2[232] <= 0;valid_bit_3[232]  <=   0;dirty_bit_3[232] <= 0;tag_address_3[232] <= 0;cache_block_3[232] <= 0;lru_counter_3[232] <= 0;valid_bit_4[232]  <=   0;dirty_bit_4[232] <= 0;tag_address_4[232] <= 0;cache_block_4[232] <= 0;lru_counter_4[232] <= 0;
        valid_bit_1[233]  <=   0;dirty_bit_1[233] <= 0;tag_address_1[233] <= 0;cache_block_1[233] <= 0;lru_counter_1[233] <= 0;valid_bit_2[233]  <=   0;dirty_bit_2[233] <= 0;tag_address_2[233] <= 0;cache_block_2[233] <= 0;lru_counter_2[233] <= 0;valid_bit_3[233]  <=   0;dirty_bit_3[233] <= 0;tag_address_3[233] <= 0;cache_block_3[233] <= 0;lru_counter_3[233] <= 0;valid_bit_4[233]  <=   0;dirty_bit_4[233] <= 0;tag_address_4[233] <= 0;cache_block_4[233] <= 0;lru_counter_4[233] <= 0;
        valid_bit_1[234]  <=   0;dirty_bit_1[234] <= 0;tag_address_1[234] <= 0;cache_block_1[234] <= 0;lru_counter_1[234] <= 0;valid_bit_2[234]  <=   0;dirty_bit_2[234] <= 0;tag_address_2[234] <= 0;cache_block_2[234] <= 0;lru_counter_2[234] <= 0;valid_bit_3[234]  <=   0;dirty_bit_3[234] <= 0;tag_address_3[234] <= 0;cache_block_3[234] <= 0;lru_counter_3[234] <= 0;valid_bit_4[234]  <=   0;dirty_bit_4[234] <= 0;tag_address_4[234] <= 0;cache_block_4[234] <= 0;lru_counter_4[234] <= 0;
        valid_bit_1[235]  <=   0;dirty_bit_1[235] <= 0;tag_address_1[235] <= 0;cache_block_1[235] <= 0;lru_counter_1[235] <= 0;valid_bit_2[235]  <=   0;dirty_bit_2[235] <= 0;tag_address_2[235] <= 0;cache_block_2[235] <= 0;lru_counter_2[235] <= 0;valid_bit_3[235]  <=   0;dirty_bit_3[235] <= 0;tag_address_3[235] <= 0;cache_block_3[235] <= 0;lru_counter_3[235] <= 0;valid_bit_4[235]  <=   0;dirty_bit_4[235] <= 0;tag_address_4[235] <= 0;cache_block_4[235] <= 0;lru_counter_4[235] <= 0;
        valid_bit_1[236]  <=   0;dirty_bit_1[236] <= 0;tag_address_1[236] <= 0;cache_block_1[236] <= 0;lru_counter_1[236] <= 0;valid_bit_2[236]  <=   0;dirty_bit_2[236] <= 0;tag_address_2[236] <= 0;cache_block_2[236] <= 0;lru_counter_2[236] <= 0;valid_bit_3[236]  <=   0;dirty_bit_3[236] <= 0;tag_address_3[236] <= 0;cache_block_3[236] <= 0;lru_counter_3[236] <= 0;valid_bit_4[236]  <=   0;dirty_bit_4[236] <= 0;tag_address_4[236] <= 0;cache_block_4[236] <= 0;lru_counter_4[236] <= 0;
        valid_bit_1[237]  <=   0;dirty_bit_1[237] <= 0;tag_address_1[237] <= 0;cache_block_1[237] <= 0;lru_counter_1[237] <= 0;valid_bit_2[237]  <=   0;dirty_bit_2[237] <= 0;tag_address_2[237] <= 0;cache_block_2[237] <= 0;lru_counter_2[237] <= 0;valid_bit_3[237]  <=   0;dirty_bit_3[237] <= 0;tag_address_3[237] <= 0;cache_block_3[237] <= 0;lru_counter_3[237] <= 0;valid_bit_4[237]  <=   0;dirty_bit_4[237] <= 0;tag_address_4[237] <= 0;cache_block_4[237] <= 0;lru_counter_4[237] <= 0;
        valid_bit_1[238]  <=   0;dirty_bit_1[238] <= 0;tag_address_1[238] <= 0;cache_block_1[238] <= 0;lru_counter_1[238] <= 0;valid_bit_2[238]  <=   0;dirty_bit_2[238] <= 0;tag_address_2[238] <= 0;cache_block_2[238] <= 0;lru_counter_2[238] <= 0;valid_bit_3[238]  <=   0;dirty_bit_3[238] <= 0;tag_address_3[238] <= 0;cache_block_3[238] <= 0;lru_counter_3[238] <= 0;valid_bit_4[238]  <=   0;dirty_bit_4[238] <= 0;tag_address_4[238] <= 0;cache_block_4[238] <= 0;lru_counter_4[238] <= 0;
        valid_bit_1[239]  <=   0;dirty_bit_1[239] <= 0;tag_address_1[239] <= 0;cache_block_1[239] <= 0;lru_counter_1[239] <= 0;valid_bit_2[239]  <=   0;dirty_bit_2[239] <= 0;tag_address_2[239] <= 0;cache_block_2[239] <= 0;lru_counter_2[239] <= 0;valid_bit_3[239]  <=   0;dirty_bit_3[239] <= 0;tag_address_3[239] <= 0;cache_block_3[239] <= 0;lru_counter_3[239] <= 0;valid_bit_4[239]  <=   0;dirty_bit_4[239] <= 0;tag_address_4[239] <= 0;cache_block_4[239] <= 0;lru_counter_4[239] <= 0;
        valid_bit_1[240]  <=   0;dirty_bit_1[240] <= 0;tag_address_1[240] <= 0;cache_block_1[240] <= 0;lru_counter_1[240] <= 0;valid_bit_2[240]  <=   0;dirty_bit_2[240] <= 0;tag_address_2[240] <= 0;cache_block_2[240] <= 0;lru_counter_2[240] <= 0;valid_bit_3[240]  <=   0;dirty_bit_3[240] <= 0;tag_address_3[240] <= 0;cache_block_3[240] <= 0;lru_counter_3[240] <= 0;valid_bit_4[240]  <=   0;dirty_bit_4[240] <= 0;tag_address_4[240] <= 0;cache_block_4[240] <= 0;lru_counter_4[240] <= 0;
        valid_bit_1[241]  <=   0;dirty_bit_1[241] <= 0;tag_address_1[241] <= 0;cache_block_1[241] <= 0;lru_counter_1[241] <= 0;valid_bit_2[241]  <=   0;dirty_bit_2[241] <= 0;tag_address_2[241] <= 0;cache_block_2[241] <= 0;lru_counter_2[241] <= 0;valid_bit_3[241]  <=   0;dirty_bit_3[241] <= 0;tag_address_3[241] <= 0;cache_block_3[241] <= 0;lru_counter_3[241] <= 0;valid_bit_4[241]  <=   0;dirty_bit_4[241] <= 0;tag_address_4[241] <= 0;cache_block_4[241] <= 0;lru_counter_4[241] <= 0;
        valid_bit_1[242]  <=   0;dirty_bit_1[242] <= 0;tag_address_1[242] <= 0;cache_block_1[242] <= 0;lru_counter_1[242] <= 0;valid_bit_2[242]  <=   0;dirty_bit_2[242] <= 0;tag_address_2[242] <= 0;cache_block_2[242] <= 0;lru_counter_2[242] <= 0;valid_bit_3[242]  <=   0;dirty_bit_3[242] <= 0;tag_address_3[242] <= 0;cache_block_3[242] <= 0;lru_counter_3[242] <= 0;valid_bit_4[242]  <=   0;dirty_bit_4[242] <= 0;tag_address_4[242] <= 0;cache_block_4[242] <= 0;lru_counter_4[242] <= 0;
        valid_bit_1[243]  <=   0;dirty_bit_1[243] <= 0;tag_address_1[243] <= 0;cache_block_1[243] <= 0;lru_counter_1[243] <= 0;valid_bit_2[243]  <=   0;dirty_bit_2[243] <= 0;tag_address_2[243] <= 0;cache_block_2[243] <= 0;lru_counter_2[243] <= 0;valid_bit_3[243]  <=   0;dirty_bit_3[243] <= 0;tag_address_3[243] <= 0;cache_block_3[243] <= 0;lru_counter_3[243] <= 0;valid_bit_4[243]  <=   0;dirty_bit_4[243] <= 0;tag_address_4[243] <= 0;cache_block_4[243] <= 0;lru_counter_4[243] <= 0;
        valid_bit_1[244]  <=   0;dirty_bit_1[244] <= 0;tag_address_1[244] <= 0;cache_block_1[244] <= 0;lru_counter_1[244] <= 0;valid_bit_2[244]  <=   0;dirty_bit_2[244] <= 0;tag_address_2[244] <= 0;cache_block_2[244] <= 0;lru_counter_2[244] <= 0;valid_bit_3[244]  <=   0;dirty_bit_3[244] <= 0;tag_address_3[244] <= 0;cache_block_3[244] <= 0;lru_counter_3[244] <= 0;valid_bit_4[244]  <=   0;dirty_bit_4[244] <= 0;tag_address_4[244] <= 0;cache_block_4[244] <= 0;lru_counter_4[244] <= 0;
        valid_bit_1[245]  <=   0;dirty_bit_1[245] <= 0;tag_address_1[245] <= 0;cache_block_1[245] <= 0;lru_counter_1[245] <= 0;valid_bit_2[245]  <=   0;dirty_bit_2[245] <= 0;tag_address_2[245] <= 0;cache_block_2[245] <= 0;lru_counter_2[245] <= 0;valid_bit_3[245]  <=   0;dirty_bit_3[245] <= 0;tag_address_3[245] <= 0;cache_block_3[245] <= 0;lru_counter_3[245] <= 0;valid_bit_4[245]  <=   0;dirty_bit_4[245] <= 0;tag_address_4[245] <= 0;cache_block_4[245] <= 0;lru_counter_4[245] <= 0;
        valid_bit_1[246]  <=   0;dirty_bit_1[246] <= 0;tag_address_1[246] <= 0;cache_block_1[246] <= 0;lru_counter_1[246] <= 0;valid_bit_2[246]  <=   0;dirty_bit_2[246] <= 0;tag_address_2[246] <= 0;cache_block_2[246] <= 0;lru_counter_2[246] <= 0;valid_bit_3[246]  <=   0;dirty_bit_3[246] <= 0;tag_address_3[246] <= 0;cache_block_3[246] <= 0;lru_counter_3[246] <= 0;valid_bit_4[246]  <=   0;dirty_bit_4[246] <= 0;tag_address_4[246] <= 0;cache_block_4[246] <= 0;lru_counter_4[246] <= 0;
        valid_bit_1[247]  <=   0;dirty_bit_1[247] <= 0;tag_address_1[247] <= 0;cache_block_1[247] <= 0;lru_counter_1[247] <= 0;valid_bit_2[247]  <=   0;dirty_bit_2[247] <= 0;tag_address_2[247] <= 0;cache_block_2[247] <= 0;lru_counter_2[247] <= 0;valid_bit_3[247]  <=   0;dirty_bit_3[247] <= 0;tag_address_3[247] <= 0;cache_block_3[247] <= 0;lru_counter_3[247] <= 0;valid_bit_4[247]  <=   0;dirty_bit_4[247] <= 0;tag_address_4[247] <= 0;cache_block_4[247] <= 0;lru_counter_4[247] <= 0;
        valid_bit_1[248]  <=   0;dirty_bit_1[248] <= 0;tag_address_1[248] <= 0;cache_block_1[248] <= 0;lru_counter_1[248] <= 0;valid_bit_2[248]  <=   0;dirty_bit_2[248] <= 0;tag_address_2[248] <= 0;cache_block_2[248] <= 0;lru_counter_2[248] <= 0;valid_bit_3[248]  <=   0;dirty_bit_3[248] <= 0;tag_address_3[248] <= 0;cache_block_3[248] <= 0;lru_counter_3[248] <= 0;valid_bit_4[248]  <=   0;dirty_bit_4[248] <= 0;tag_address_4[248] <= 0;cache_block_4[248] <= 0;lru_counter_4[248] <= 0;
        valid_bit_1[249]  <=   0;dirty_bit_1[249] <= 0;tag_address_1[249] <= 0;cache_block_1[249] <= 0;lru_counter_1[249] <= 0;valid_bit_2[249]  <=   0;dirty_bit_2[249] <= 0;tag_address_2[249] <= 0;cache_block_2[249] <= 0;lru_counter_2[249] <= 0;valid_bit_3[249]  <=   0;dirty_bit_3[249] <= 0;tag_address_3[249] <= 0;cache_block_3[249] <= 0;lru_counter_3[249] <= 0;valid_bit_4[249]  <=   0;dirty_bit_4[249] <= 0;tag_address_4[249] <= 0;cache_block_4[249] <= 0;lru_counter_4[249] <= 0;
        valid_bit_1[250]  <=   0;dirty_bit_1[250] <= 0;tag_address_1[250] <= 0;cache_block_1[250] <= 0;lru_counter_1[250] <= 0;valid_bit_2[250]  <=   0;dirty_bit_2[250] <= 0;tag_address_2[250] <= 0;cache_block_2[250] <= 0;lru_counter_2[250] <= 0;valid_bit_3[250]  <=   0;dirty_bit_3[250] <= 0;tag_address_3[250] <= 0;cache_block_3[250] <= 0;lru_counter_3[250] <= 0;valid_bit_4[250]  <=   0;dirty_bit_4[250] <= 0;tag_address_4[250] <= 0;cache_block_4[250] <= 0;lru_counter_4[250] <= 0;
        valid_bit_1[251]  <=   0;dirty_bit_1[251] <= 0;tag_address_1[251] <= 0;cache_block_1[251] <= 0;lru_counter_1[251] <= 0;valid_bit_2[251]  <=   0;dirty_bit_2[251] <= 0;tag_address_2[251] <= 0;cache_block_2[251] <= 0;lru_counter_2[251] <= 0;valid_bit_3[251]  <=   0;dirty_bit_3[251] <= 0;tag_address_3[251] <= 0;cache_block_3[251] <= 0;lru_counter_3[251] <= 0;valid_bit_4[251]  <=   0;dirty_bit_4[251] <= 0;tag_address_4[251] <= 0;cache_block_4[251] <= 0;lru_counter_4[251] <= 0;
        valid_bit_1[252]  <=   0;dirty_bit_1[252] <= 0;tag_address_1[252] <= 0;cache_block_1[252] <= 0;lru_counter_1[252] <= 0;valid_bit_2[252]  <=   0;dirty_bit_2[252] <= 0;tag_address_2[252] <= 0;cache_block_2[252] <= 0;lru_counter_2[252] <= 0;valid_bit_3[252]  <=   0;dirty_bit_3[252] <= 0;tag_address_3[252] <= 0;cache_block_3[252] <= 0;lru_counter_3[252] <= 0;valid_bit_4[252]  <=   0;dirty_bit_4[252] <= 0;tag_address_4[252] <= 0;cache_block_4[252] <= 0;lru_counter_4[252] <= 0;
        valid_bit_1[253]  <=   0;dirty_bit_1[253] <= 0;tag_address_1[253] <= 0;cache_block_1[253] <= 0;lru_counter_1[253] <= 0;valid_bit_2[253]  <=   0;dirty_bit_2[253] <= 0;tag_address_2[253] <= 0;cache_block_2[253] <= 0;lru_counter_2[253] <= 0;valid_bit_3[253]  <=   0;dirty_bit_3[253] <= 0;tag_address_3[253] <= 0;cache_block_3[253] <= 0;lru_counter_3[253] <= 0;valid_bit_4[253]  <=   0;dirty_bit_4[253] <= 0;tag_address_4[253] <= 0;cache_block_4[253] <= 0;lru_counter_4[253] <= 0;
        valid_bit_1[254]  <=   0;dirty_bit_1[254] <= 0;tag_address_1[254] <= 0;cache_block_1[254] <= 0;lru_counter_1[254] <= 0;valid_bit_2[254]  <=   0;dirty_bit_2[254] <= 0;tag_address_2[254] <= 0;cache_block_2[254] <= 0;lru_counter_2[254] <= 0;valid_bit_3[254]  <=   0;dirty_bit_3[254] <= 0;tag_address_3[254] <= 0;cache_block_3[254] <= 0;lru_counter_3[254] <= 0;valid_bit_4[254]  <=   0;dirty_bit_4[254] <= 0;tag_address_4[254] <= 0;cache_block_4[254] <= 0;lru_counter_4[254] <= 0;
        valid_bit_1[255]  <=   0;dirty_bit_1[255] <= 0;tag_address_1[255] <= 0;cache_block_1[255] <= 0;lru_counter_1[255] <= 0;valid_bit_2[255]  <=   0;dirty_bit_2[255] <= 0;tag_address_2[255] <= 0;cache_block_2[255] <= 0;lru_counter_2[255] <= 0;valid_bit_3[255]  <=   0;dirty_bit_3[255] <= 0;tag_address_3[255] <= 0;cache_block_3[255] <= 0;lru_counter_3[255] <= 0;valid_bit_4[255]  <=   0;dirty_bit_4[255] <= 0;tag_address_4[255] <= 0;cache_block_4[255] <= 0;lru_counter_4[255] <= 0;
    end
end


endmodule


/*
else begin
    //wr miss
    //wr allocate
    if(!valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
        //block 1
        cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        valid_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        o_mem_wr_en                                                            <=   0;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2; 
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1;
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0; 
    end
    else if(!valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
        cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        valid_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        o_mem_wr_en                                                            <=   0;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2;
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3; 
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1;
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0; 
    end
    else if(!valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
        cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        valid_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        o_mem_wr_en                                                            <=   0;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1;
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2; 
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0; 
    end
    else if(!valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
        cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        valid_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        o_mem_wr_en                                                            <=   0;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 0;
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 1; 
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 2;
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3; 
    end
    else if(lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
        if(dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
            o_mem_wr_data <= cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
            o_mem_wr_address <= {tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
            o_mem_wr_en <= 1;
        end
        cache_block_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
    
    end
    else if(lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
        if(dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
            o_mem_wr_data <= cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
            o_mem_wr_address <= {tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
            o_mem_wr_en <= 1;
        end
        cache_block_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
    end
    else if(lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
        if(dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
            o_mem_wr_data <= cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
            o_mem_wr_address <= {tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
            o_mem_wr_en <= 1;
        end
        cache_block_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
    end
    else if(lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]==0) begin
        if(dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]) begin
            o_mem_wr_data <= cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
            o_mem_wr_address <= {tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]],i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW],6'd0};
            o_mem_wr_en <= 1;
        end
        cache_block_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_wr_data;
        tag_address_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]       <=   i_cpu_address[TAG_HIGH:TAG_LOW];
        dirty_bit_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]         <=   1;
        o_cpu_busy                                                             <=   0;
        lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= 3;
        lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_1[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_2[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
        lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]]  <= (lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] > lru_counter_4[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]])? lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]] -1 : lru_counter_3[i_cpu_address[BLOCK_ADDRESS_HIGH:BLOCK_ADDRESS_LOW]];
    end
end

*/
